module NV_NVDLA_SDP_CORE_Y_lut(nvdla_core_clk, nvdla_core_rstn, idx2lut_pd, idx2lut_pvld, lut2inp_prdy, op_en_load, pwrbus_ram_pd, reg2dp_lut_int_access_type, reg2dp_lut_int_addr, reg2dp_lut_int_data, reg2dp_lut_int_data_wr, reg2dp_lut_int_table_id, reg2dp_lut_le_end, reg2dp_lut_le_function, reg2dp_lut_le_index_offset, reg2dp_lut_le_slope_oflow_scale, reg2dp_lut_le_slope_oflow_shift, reg2dp_lut_le_slope_uflow_scale, reg2dp_lut_le_slope_uflow_shift, reg2dp_lut_le_start, reg2dp_lut_lo_end, reg2dp_lut_lo_slope_oflow_scale, reg2dp_lut_lo_slope_oflow_shift, reg2dp_lut_lo_slope_uflow_scale, reg2dp_lut_lo_slope_uflow_shift, reg2dp_lut_lo_start, reg2dp_perf_lut_en, reg2dp_proc_precision, dp2reg_lut_hybrid, dp2reg_lut_int_data, dp2reg_lut_le_hit, dp2reg_lut_lo_hit, dp2reg_lut_oflow, dp2reg_lut_uflow, idx2lut_prdy, lut2inp_pd, lut2inp_pvld);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1867" *)
  wire [15:0] _0000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2487" *)
  wire [15:0] _0001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2549" *)
  wire [15:0] _0002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2611" *)
  wire [15:0] _0003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2673" *)
  wire [15:0] _0004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2735" *)
  wire [15:0] _0005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2797" *)
  wire [15:0] _0006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2859" *)
  wire [15:0] _0007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2921" *)
  wire [15:0] _0008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2983" *)
  wire [15:0] _0009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3045" *)
  wire [15:0] _0010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1929" *)
  wire [15:0] _0011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3107" *)
  wire [15:0] _0012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3169" *)
  wire [15:0] _0013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3231" *)
  wire [15:0] _0014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3293" *)
  wire [15:0] _0015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3355" *)
  wire [15:0] _0016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3417" *)
  wire [15:0] _0017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3479" *)
  wire [15:0] _0018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3541" *)
  wire [15:0] _0019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3603" *)
  wire [15:0] _0020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3665" *)
  wire [15:0] _0021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1991" *)
  wire [15:0] _0022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3727" *)
  wire [15:0] _0023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3789" *)
  wire [15:0] _0024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3851" *)
  wire [15:0] _0025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3913" *)
  wire [15:0] _0026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3975" *)
  wire [15:0] _0027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4037" *)
  wire [15:0] _0028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4099" *)
  wire [15:0] _0029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4161" *)
  wire [15:0] _0030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4223" *)
  wire [15:0] _0031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4285" *)
  wire [15:0] _0032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2053" *)
  wire [15:0] _0033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4347" *)
  wire [15:0] _0034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4409" *)
  wire [15:0] _0035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4471" *)
  wire [15:0] _0036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4533" *)
  wire [15:0] _0037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4595" *)
  wire [15:0] _0038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4657" *)
  wire [15:0] _0039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4719" *)
  wire [15:0] _0040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4781" *)
  wire [15:0] _0041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4843" *)
  wire [15:0] _0042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4905" *)
  wire [15:0] _0043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2115" *)
  wire [15:0] _0044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4967" *)
  wire [15:0] _0045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5029" *)
  wire [15:0] _0046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5091" *)
  wire [15:0] _0047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5153" *)
  wire [15:0] _0048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5215" *)
  wire [15:0] _0049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5277" *)
  wire [15:0] _0050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5339" *)
  wire [15:0] _0051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5401" *)
  wire [15:0] _0052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5463" *)
  wire [15:0] _0053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5525" *)
  wire [15:0] _0054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2177" *)
  wire [15:0] _0055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5587" *)
  wire [15:0] _0056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5649" *)
  wire [15:0] _0057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5711" *)
  wire [15:0] _0058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5773" *)
  wire [15:0] _0059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5835" *)
  wire [15:0] _0060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2239" *)
  wire [15:0] _0061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2301" *)
  wire [15:0] _0062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2363" *)
  wire [15:0] _0063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2425" *)
  wire [15:0] _0064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6089" *)
  wire [15:0] _0065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12289" *)
  wire [15:0] _0066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12351" *)
  wire [15:0] _0067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12413" *)
  wire [15:0] _0068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12475" *)
  wire [15:0] _0069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12537" *)
  wire [15:0] _0070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12599" *)
  wire [15:0] _0071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12661" *)
  wire [15:0] _0072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12723" *)
  wire [15:0] _0073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12785" *)
  wire [15:0] _0074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12847" *)
  wire [15:0] _0075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6709" *)
  wire [15:0] _0076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12909" *)
  wire [15:0] _0077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12971" *)
  wire [15:0] _0078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13033" *)
  wire [15:0] _0079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13095" *)
  wire [15:0] _0080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13157" *)
  wire [15:0] _0081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13219" *)
  wire [15:0] _0082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13281" *)
  wire [15:0] _0083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13343" *)
  wire [15:0] _0084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13405" *)
  wire [15:0] _0085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13467" *)
  wire [15:0] _0086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6771" *)
  wire [15:0] _0087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13529" *)
  wire [15:0] _0088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13591" *)
  wire [15:0] _0089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13653" *)
  wire [15:0] _0090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13715" *)
  wire [15:0] _0091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13777" *)
  wire [15:0] _0092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13839" *)
  wire [15:0] _0093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13901" *)
  wire [15:0] _0094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13963" *)
  wire [15:0] _0095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14025" *)
  wire [15:0] _0096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14087" *)
  wire [15:0] _0097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6833" *)
  wire [15:0] _0098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14149" *)
  wire [15:0] _0099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14211" *)
  wire [15:0] _0100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14273" *)
  wire [15:0] _0101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14335" *)
  wire [15:0] _0102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14397" *)
  wire [15:0] _0103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14459" *)
  wire [15:0] _0104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14521" *)
  wire [15:0] _0105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14583" *)
  wire [15:0] _0106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14645" *)
  wire [15:0] _0107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14707" *)
  wire [15:0] _0108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6895" *)
  wire [15:0] _0109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14769" *)
  wire [15:0] _0110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14831" *)
  wire [15:0] _0111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14893" *)
  wire [15:0] _0112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14955" *)
  wire [15:0] _0113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15017" *)
  wire [15:0] _0114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15079" *)
  wire [15:0] _0115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15141" *)
  wire [15:0] _0116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15203" *)
  wire [15:0] _0117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15265" *)
  wire [15:0] _0118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15327" *)
  wire [15:0] _0119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6957" *)
  wire [15:0] _0120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15389" *)
  wire [15:0] _0121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15451" *)
  wire [15:0] _0122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15513" *)
  wire [15:0] _0123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15575" *)
  wire [15:0] _0124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15637" *)
  wire [15:0] _0125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15699" *)
  wire [15:0] _0126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15761" *)
  wire [15:0] _0127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15823" *)
  wire [15:0] _0128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15885" *)
  wire [15:0] _0129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15947" *)
  wire [15:0] _0130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7019" *)
  wire [15:0] _0131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16009" *)
  wire [15:0] _0132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16071" *)
  wire [15:0] _0133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16133" *)
  wire [15:0] _0134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16195" *)
  wire [15:0] _0135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16257" *)
  wire [15:0] _0136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16319" *)
  wire [15:0] _0137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16381" *)
  wire [15:0] _0138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16443" *)
  wire [15:0] _0139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16505" *)
  wire [15:0] _0140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16567" *)
  wire [15:0] _0141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7081" *)
  wire [15:0] _0142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16629" *)
  wire [15:0] _0143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16691" *)
  wire [15:0] _0144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16753" *)
  wire [15:0] _0145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16815" *)
  wire [15:0] _0146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16877" *)
  wire [15:0] _0147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16939" *)
  wire [15:0] _0148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17001" *)
  wire [15:0] _0149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17063" *)
  wire [15:0] _0150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17125" *)
  wire [15:0] _0151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17187" *)
  wire [15:0] _0152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7143" *)
  wire [15:0] _0153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17249" *)
  wire [15:0] _0154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17311" *)
  wire [15:0] _0155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17373" *)
  wire [15:0] _0156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17435" *)
  wire [15:0] _0157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17497" *)
  wire [15:0] _0158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17559" *)
  wire [15:0] _0159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17621" *)
  wire [15:0] _0160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17683" *)
  wire [15:0] _0161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17745" *)
  wire [15:0] _0162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17807" *)
  wire [15:0] _0163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7205" *)
  wire [15:0] _0164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17869" *)
  wire [15:0] _0165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17931" *)
  wire [15:0] _0166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17993" *)
  wire [15:0] _0167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18055" *)
  wire [15:0] _0168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18117" *)
  wire [15:0] _0169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18179" *)
  wire [15:0] _0170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18241" *)
  wire [15:0] _0171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18303" *)
  wire [15:0] _0172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18365" *)
  wire [15:0] _0173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18427" *)
  wire [15:0] _0174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7267" *)
  wire [15:0] _0175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6151" *)
  wire [15:0] _0176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18489" *)
  wire [15:0] _0177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18551" *)
  wire [15:0] _0178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18613" *)
  wire [15:0] _0179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18675" *)
  wire [15:0] _0180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18737" *)
  wire [15:0] _0181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18799" *)
  wire [15:0] _0182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18861" *)
  wire [15:0] _0183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18923" *)
  wire [15:0] _0184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18985" *)
  wire [15:0] _0185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19047" *)
  wire [15:0] _0186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7329" *)
  wire [15:0] _0187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19109" *)
  wire [15:0] _0188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19171" *)
  wire [15:0] _0189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19233" *)
  wire [15:0] _0190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19295" *)
  wire [15:0] _0191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19357" *)
  wire [15:0] _0192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19419" *)
  wire [15:0] _0193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19481" *)
  wire [15:0] _0194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19543" *)
  wire [15:0] _0195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19605" *)
  wire [15:0] _0196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19667" *)
  wire [15:0] _0197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7391" *)
  wire [15:0] _0198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19729" *)
  wire [15:0] _0199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19791" *)
  wire [15:0] _0200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19853" *)
  wire [15:0] _0201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19915" *)
  wire [15:0] _0202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19977" *)
  wire [15:0] _0203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20039" *)
  wire [15:0] _0204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20101" *)
  wire [15:0] _0205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20163" *)
  wire [15:0] _0206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20225" *)
  wire [15:0] _0207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20287" *)
  wire [15:0] _0208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7453" *)
  wire [15:0] _0209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20349" *)
  wire [15:0] _0210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20411" *)
  wire [15:0] _0211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20473" *)
  wire [15:0] _0212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20535" *)
  wire [15:0] _0213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20597" *)
  wire [15:0] _0214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20659" *)
  wire [15:0] _0215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20721" *)
  wire [15:0] _0216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20783" *)
  wire [15:0] _0217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20845" *)
  wire [15:0] _0218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20907" *)
  wire [15:0] _0219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7515" *)
  wire [15:0] _0220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20969" *)
  wire [15:0] _0221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21031" *)
  wire [15:0] _0222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21093" *)
  wire [15:0] _0223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21155" *)
  wire [15:0] _0224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21217" *)
  wire [15:0] _0225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21279" *)
  wire [15:0] _0226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21341" *)
  wire [15:0] _0227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21403" *)
  wire [15:0] _0228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21465" *)
  wire [15:0] _0229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21527" *)
  wire [15:0] _0230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7577" *)
  wire [15:0] _0231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21589" *)
  wire [15:0] _0232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21651" *)
  wire [15:0] _0233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21713" *)
  wire [15:0] _0234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21775" *)
  wire [15:0] _0235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21837" *)
  wire [15:0] _0236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21899" *)
  wire [15:0] _0237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21961" *)
  wire [15:0] _0238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7639" *)
  wire [15:0] _0239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7701" *)
  wire [15:0] _0240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7763" *)
  wire [15:0] _0241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7825" *)
  wire [15:0] _0242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7887" *)
  wire [15:0] _0243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6213" *)
  wire [15:0] _0244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7949" *)
  wire [15:0] _0245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8011" *)
  wire [15:0] _0246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8073" *)
  wire [15:0] _0247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8135" *)
  wire [15:0] _0248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8197" *)
  wire [15:0] _0249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8259" *)
  wire [15:0] _0250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8321" *)
  wire [15:0] _0251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8383" *)
  wire [15:0] _0252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8445" *)
  wire [15:0] _0253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8507" *)
  wire [15:0] _0254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6275" *)
  wire [15:0] _0255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8569" *)
  wire [15:0] _0256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8631" *)
  wire [15:0] _0257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8693" *)
  wire [15:0] _0258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8755" *)
  wire [15:0] _0259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8817" *)
  wire [15:0] _0260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8879" *)
  wire [15:0] _0261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8941" *)
  wire [15:0] _0262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9003" *)
  wire [15:0] _0263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9065" *)
  wire [15:0] _0264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9127" *)
  wire [15:0] _0265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6337" *)
  wire [15:0] _0266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9189" *)
  wire [15:0] _0267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9251" *)
  wire [15:0] _0268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9313" *)
  wire [15:0] _0269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9375" *)
  wire [15:0] _0270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9437" *)
  wire [15:0] _0271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9499" *)
  wire [15:0] _0272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9561" *)
  wire [15:0] _0273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9623" *)
  wire [15:0] _0274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9685" *)
  wire [15:0] _0275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9747" *)
  wire [15:0] _0276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6399" *)
  wire [15:0] _0277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9809" *)
  wire [15:0] _0278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9871" *)
  wire [15:0] _0279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9933" *)
  wire [15:0] _0280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9995" *)
  wire [15:0] _0281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10057" *)
  wire [15:0] _0282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10119" *)
  wire [15:0] _0283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10181" *)
  wire [15:0] _0284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10243" *)
  wire [15:0] _0285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10305" *)
  wire [15:0] _0286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10367" *)
  wire [15:0] _0287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6461" *)
  wire [15:0] _0288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10429" *)
  wire [15:0] _0289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10491" *)
  wire [15:0] _0290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10553" *)
  wire [15:0] _0291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10615" *)
  wire [15:0] _0292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10677" *)
  wire [15:0] _0293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10739" *)
  wire [15:0] _0294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10801" *)
  wire [15:0] _0295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10863" *)
  wire [15:0] _0296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10925" *)
  wire [15:0] _0297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10987" *)
  wire [15:0] _0298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6523" *)
  wire [15:0] _0299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11049" *)
  wire [15:0] _0300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11111" *)
  wire [15:0] _0301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11173" *)
  wire [15:0] _0302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11235" *)
  wire [15:0] _0303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11297" *)
  wire [15:0] _0304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11359" *)
  wire [15:0] _0305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11421" *)
  wire [15:0] _0306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11483" *)
  wire [15:0] _0307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11545" *)
  wire [15:0] _0308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11607" *)
  wire [15:0] _0309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6585" *)
  wire [15:0] _0310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11669" *)
  wire [15:0] _0311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11731" *)
  wire [15:0] _0312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11793" *)
  wire [15:0] _0313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11855" *)
  wire [15:0] _0314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11917" *)
  wire [15:0] _0315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11979" *)
  wire [15:0] _0316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12041" *)
  wire [15:0] _0317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12103" *)
  wire [15:0] _0318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12165" *)
  wire [15:0] _0319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12227" *)
  wire [15:0] _0320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6647" *)
  wire [15:0] _0321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [7:0] _0322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22228" *)
  wire [323:0] _0323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22221" *)
  wire _0324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31592" *)
  wire [739:0] _0325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31585" *)
  wire _0326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31623" *)
  wire [739:0] _0327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31612" *)
  wire _0328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22497" *)
  wire [31:0] _0329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22540" *)
  wire [31:0] _0330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22583" *)
  wire [31:0] _0331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22407" *)
  wire [31:0] _0332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22450" *)
  wire [31:0] _0333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [31:0] _0335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [31:0] _0336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [31:0] _0337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [31:0] _0339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [31:0] _0340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [31:0] _0341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [15:0] _0342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [15:0] _0343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [15:0] _0344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [15:0] _0345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [4:0] _0346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [4:0] _0347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [4:0] _0348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [4:0] _0349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [31:0] _0352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [31:0] _0353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [31:0] _0354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [15:0] _0355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [15:0] _0356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [15:0] _0357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [15:0] _0358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [4:0] _0359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [4:0] _0360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [4:0] _0361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [4:0] _0362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [31:0] _0364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [31:0] _0365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [31:0] _0366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [31:0] _0367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [15:0] _0368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [15:0] _0369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [15:0] _0370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [15:0] _0371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31100" *)
  wire [4:0] _0372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31162" *)
  wire [4:0] _0373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31224" *)
  wire [4:0] _0374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31286" *)
  wire [4:0] _0375_;
  wire [1:0] _0376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22380" *)
  wire [2:0] _0377_;
  wire [1:0] _0378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22423" *)
  wire [2:0] _0379_;
  wire [1:0] _0380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22470" *)
  wire [2:0] _0381_;
  wire [1:0] _0382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22513" *)
  wire [2:0] _0383_;
  wire [1:0] _0384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22556" *)
  wire [2:0] _0385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10056" *)
  wire _0386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1866" *)
  wire _0387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10056" *)
  wire _0388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10118" *)
  wire _0389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10180" *)
  wire _0390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10242" *)
  wire _0391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10304" *)
  wire _0392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10366" *)
  wire _0393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10428" *)
  wire _0394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10490" *)
  wire _0395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10552" *)
  wire _0396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10614" *)
  wire _0397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10676" *)
  wire _0398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10738" *)
  wire _0399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10800" *)
  wire _0400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10862" *)
  wire _0401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10924" *)
  wire _0402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10986" *)
  wire _0403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11048" *)
  wire _0404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11110" *)
  wire _0405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11172" *)
  wire _0406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11234" *)
  wire _0407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11296" *)
  wire _0408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11358" *)
  wire _0409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11420" *)
  wire _0410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11482" *)
  wire _0411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11544" *)
  wire _0412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11606" *)
  wire _0413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11668" *)
  wire _0414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11730" *)
  wire _0415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11792" *)
  wire _0416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11854" *)
  wire _0417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11916" *)
  wire _0418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11978" *)
  wire _0419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12040" *)
  wire _0420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12102" *)
  wire _0421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12164" *)
  wire _0422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12226" *)
  wire _0423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12288" *)
  wire _0424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12350" *)
  wire _0425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12412" *)
  wire _0426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12474" *)
  wire _0427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12536" *)
  wire _0428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12598" *)
  wire _0429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12660" *)
  wire _0430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12722" *)
  wire _0431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12784" *)
  wire _0432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12846" *)
  wire _0433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12908" *)
  wire _0434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12970" *)
  wire _0435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13032" *)
  wire _0436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13094" *)
  wire _0437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13156" *)
  wire _0438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13218" *)
  wire _0439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13280" *)
  wire _0440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13342" *)
  wire _0441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13404" *)
  wire _0442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13466" *)
  wire _0443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13528" *)
  wire _0444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13590" *)
  wire _0445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13652" *)
  wire _0446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13714" *)
  wire _0447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13776" *)
  wire _0448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13838" *)
  wire _0449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13900" *)
  wire _0450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13962" *)
  wire _0451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14024" *)
  wire _0452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14086" *)
  wire _0453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14148" *)
  wire _0454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14210" *)
  wire _0455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14272" *)
  wire _0456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14334" *)
  wire _0457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14396" *)
  wire _0458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14458" *)
  wire _0459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14520" *)
  wire _0460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14582" *)
  wire _0461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14644" *)
  wire _0462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14706" *)
  wire _0463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14768" *)
  wire _0464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14830" *)
  wire _0465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14892" *)
  wire _0466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14954" *)
  wire _0467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15016" *)
  wire _0468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15078" *)
  wire _0469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15140" *)
  wire _0470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15202" *)
  wire _0471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15264" *)
  wire _0472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15326" *)
  wire _0473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15388" *)
  wire _0474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15450" *)
  wire _0475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15512" *)
  wire _0476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15574" *)
  wire _0477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15636" *)
  wire _0478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15698" *)
  wire _0479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15760" *)
  wire _0480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15822" *)
  wire _0481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15884" *)
  wire _0482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15946" *)
  wire _0483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16008" *)
  wire _0484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16070" *)
  wire _0485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16132" *)
  wire _0486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16194" *)
  wire _0487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16256" *)
  wire _0488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16318" *)
  wire _0489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16380" *)
  wire _0490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16442" *)
  wire _0491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16504" *)
  wire _0492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16566" *)
  wire _0493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16628" *)
  wire _0494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16690" *)
  wire _0495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16752" *)
  wire _0496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16814" *)
  wire _0497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16876" *)
  wire _0498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16938" *)
  wire _0499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17000" *)
  wire _0500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17062" *)
  wire _0501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17124" *)
  wire _0502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17186" *)
  wire _0503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17248" *)
  wire _0504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17310" *)
  wire _0505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17372" *)
  wire _0506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17434" *)
  wire _0507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17496" *)
  wire _0508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17558" *)
  wire _0509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17620" *)
  wire _0510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17682" *)
  wire _0511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17744" *)
  wire _0512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17806" *)
  wire _0513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17868" *)
  wire _0514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17930" *)
  wire _0515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17992" *)
  wire _0516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18054" *)
  wire _0517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18116" *)
  wire _0518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18178" *)
  wire _0519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18240" *)
  wire _0520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18302" *)
  wire _0521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18364" *)
  wire _0522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18426" *)
  wire _0523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18488" *)
  wire _0524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18550" *)
  wire _0525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18612" *)
  wire _0526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1866" *)
  wire _0527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18674" *)
  wire _0528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18736" *)
  wire _0529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18798" *)
  wire _0530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18860" *)
  wire _0531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18922" *)
  wire _0532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18984" *)
  wire _0533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19046" *)
  wire _0534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19108" *)
  wire _0535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19170" *)
  wire _0536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19232" *)
  wire _0537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1928" *)
  wire _0538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19294" *)
  wire _0539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19356" *)
  wire _0540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19418" *)
  wire _0541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19480" *)
  wire _0542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19542" *)
  wire _0543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19604" *)
  wire _0544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19666" *)
  wire _0545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19728" *)
  wire _0546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19790" *)
  wire _0547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19852" *)
  wire _0548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1990" *)
  wire _0549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19914" *)
  wire _0550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19976" *)
  wire _0551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20038" *)
  wire _0552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20100" *)
  wire _0553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20162" *)
  wire _0554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20224" *)
  wire _0555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20286" *)
  wire _0556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20348" *)
  wire _0557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20410" *)
  wire _0558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20472" *)
  wire _0559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2052" *)
  wire _0560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20534" *)
  wire _0561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20596" *)
  wire _0562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20658" *)
  wire _0563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20720" *)
  wire _0564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20782" *)
  wire _0565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20844" *)
  wire _0566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20906" *)
  wire _0567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20968" *)
  wire _0568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21030" *)
  wire _0569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21092" *)
  wire _0570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2114" *)
  wire _0571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21154" *)
  wire _0572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21216" *)
  wire _0573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21278" *)
  wire _0574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21340" *)
  wire _0575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21402" *)
  wire _0576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21464" *)
  wire _0577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21526" *)
  wire _0578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21588" *)
  wire _0579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21650" *)
  wire _0580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21712" *)
  wire _0581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2176" *)
  wire _0582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21774" *)
  wire _0583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21836" *)
  wire _0584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21898" *)
  wire _0585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21960" *)
  wire _0586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2238" *)
  wire _0587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2300" *)
  wire _0588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2362" *)
  wire _0589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2424" *)
  wire _0590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2486" *)
  wire _0591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2548" *)
  wire _0592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2610" *)
  wire _0593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2672" *)
  wire _0594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2734" *)
  wire _0595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2796" *)
  wire _0596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2858" *)
  wire _0597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2920" *)
  wire _0598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2982" *)
  wire _0599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3044" *)
  wire _0600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3106" *)
  wire _0601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31126" *)
  wire _0602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3168" *)
  wire _0603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3230" *)
  wire _0604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3292" *)
  wire _0605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3354" *)
  wire _0606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3416" *)
  wire _0607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3478" *)
  wire _0608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3540" *)
  wire _0609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3602" *)
  wire _0610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3664" *)
  wire _0611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3726" *)
  wire _0612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3788" *)
  wire _0613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3850" *)
  wire _0614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3912" *)
  wire _0615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3974" *)
  wire _0616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4036" *)
  wire _0617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4098" *)
  wire _0618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4160" *)
  wire _0619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4222" *)
  wire _0620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4284" *)
  wire _0621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4346" *)
  wire _0622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4408" *)
  wire _0623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4470" *)
  wire _0624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4532" *)
  wire _0625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4594" *)
  wire _0626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4656" *)
  wire _0627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4718" *)
  wire _0628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4780" *)
  wire _0629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4842" *)
  wire _0630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4904" *)
  wire _0631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4966" *)
  wire _0632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5028" *)
  wire _0633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5090" *)
  wire _0634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5152" *)
  wire _0635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5214" *)
  wire _0636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5276" *)
  wire _0637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5338" *)
  wire _0638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5400" *)
  wire _0639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5462" *)
  wire _0640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5524" *)
  wire _0641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5586" *)
  wire _0642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5648" *)
  wire _0643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5710" *)
  wire _0644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5772" *)
  wire _0645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22230" *)
  wire _0646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31594" *)
  wire _0647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31609" *)
  wire _0648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22219" *)
  wire _0649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31583" *)
  wire _0650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31609" *)
  wire _0651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31610" *)
  wire _0652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22466" *)
  wire _0653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22467" *)
  wire _0654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22468" *)
  wire _0655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22469" *)
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22381" *)
  wire _2709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22424" *)
  wire _2710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22471" *)
  wire _2711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22514" *)
  wire _2712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22557" *)
  wire _2713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31132" *)
  wire [31:0] _2714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31132" *)
  wire [31:0] _2715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:89" *)
  reg [15:0] REG_le_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:90" *)
  reg [15:0] REG_le_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:91" *)
  reg [15:0] REG_le_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:520" *)
  wire [15:0] REG_le_100;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:521" *)
  wire [15:0] REG_le_101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:522" *)
  wire [15:0] REG_le_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:523" *)
  wire [15:0] REG_le_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:524" *)
  wire [15:0] REG_le_104;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:525" *)
  wire [15:0] REG_le_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:526" *)
  wire [15:0] REG_le_106;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:527" *)
  wire [15:0] REG_le_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:528" *)
  wire [15:0] REG_le_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:529" *)
  wire [15:0] REG_le_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:92" *)
  reg [15:0] REG_le_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:530" *)
  wire [15:0] REG_le_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:531" *)
  wire [15:0] REG_le_111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:532" *)
  wire [15:0] REG_le_112;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:533" *)
  wire [15:0] REG_le_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:534" *)
  wire [15:0] REG_le_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:535" *)
  wire [15:0] REG_le_115;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:536" *)
  wire [15:0] REG_le_116;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:537" *)
  wire [15:0] REG_le_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:538" *)
  wire [15:0] REG_le_118;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:539" *)
  wire [15:0] REG_le_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:93" *)
  reg [15:0] REG_le_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:540" *)
  wire [15:0] REG_le_120;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:541" *)
  wire [15:0] REG_le_121;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:542" *)
  wire [15:0] REG_le_122;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:543" *)
  wire [15:0] REG_le_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:544" *)
  wire [15:0] REG_le_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:545" *)
  wire [15:0] REG_le_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:546" *)
  wire [15:0] REG_le_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:547" *)
  wire [15:0] REG_le_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:548" *)
  wire [15:0] REG_le_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:549" *)
  wire [15:0] REG_le_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:94" *)
  reg [15:0] REG_le_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:550" *)
  wire [15:0] REG_le_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:551" *)
  wire [15:0] REG_le_131;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:552" *)
  wire [15:0] REG_le_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:553" *)
  wire [15:0] REG_le_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:554" *)
  wire [15:0] REG_le_134;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:555" *)
  wire [15:0] REG_le_135;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:556" *)
  wire [15:0] REG_le_136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:557" *)
  wire [15:0] REG_le_137;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:558" *)
  wire [15:0] REG_le_138;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:559" *)
  wire [15:0] REG_le_139;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:95" *)
  reg [15:0] REG_le_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:560" *)
  wire [15:0] REG_le_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:561" *)
  wire [15:0] REG_le_141;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:562" *)
  wire [15:0] REG_le_142;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:563" *)
  wire [15:0] REG_le_143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:564" *)
  wire [15:0] REG_le_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:565" *)
  wire [15:0] REG_le_145;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:566" *)
  wire [15:0] REG_le_146;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:567" *)
  wire [15:0] REG_le_147;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:568" *)
  wire [15:0] REG_le_148;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:569" *)
  wire [15:0] REG_le_149;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:96" *)
  reg [15:0] REG_le_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:570" *)
  wire [15:0] REG_le_150;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:571" *)
  wire [15:0] REG_le_151;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:572" *)
  wire [15:0] REG_le_152;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:573" *)
  wire [15:0] REG_le_153;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:574" *)
  wire [15:0] REG_le_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:575" *)
  wire [15:0] REG_le_155;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:576" *)
  wire [15:0] REG_le_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:577" *)
  wire [15:0] REG_le_157;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:578" *)
  wire [15:0] REG_le_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:579" *)
  wire [15:0] REG_le_159;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:97" *)
  reg [15:0] REG_le_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:580" *)
  wire [15:0] REG_le_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:581" *)
  wire [15:0] REG_le_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:582" *)
  wire [15:0] REG_le_162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:583" *)
  wire [15:0] REG_le_163;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:584" *)
  wire [15:0] REG_le_164;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:585" *)
  wire [15:0] REG_le_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:586" *)
  wire [15:0] REG_le_166;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:587" *)
  wire [15:0] REG_le_167;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:588" *)
  wire [15:0] REG_le_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:589" *)
  wire [15:0] REG_le_169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:98" *)
  reg [15:0] REG_le_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:590" *)
  wire [15:0] REG_le_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:591" *)
  wire [15:0] REG_le_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:592" *)
  wire [15:0] REG_le_172;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:593" *)
  wire [15:0] REG_le_173;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:594" *)
  wire [15:0] REG_le_174;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:595" *)
  wire [15:0] REG_le_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:596" *)
  wire [15:0] REG_le_176;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:597" *)
  wire [15:0] REG_le_177;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:598" *)
  wire [15:0] REG_le_178;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:599" *)
  wire [15:0] REG_le_179;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:99" *)
  reg [15:0] REG_le_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:600" *)
  wire [15:0] REG_le_180;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:601" *)
  wire [15:0] REG_le_181;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:602" *)
  wire [15:0] REG_le_182;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:603" *)
  wire [15:0] REG_le_183;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:604" *)
  wire [15:0] REG_le_184;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:605" *)
  wire [15:0] REG_le_185;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:606" *)
  wire [15:0] REG_le_186;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:607" *)
  wire [15:0] REG_le_187;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:608" *)
  wire [15:0] REG_le_188;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:609" *)
  wire [15:0] REG_le_189;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:100" *)
  reg [15:0] REG_le_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:610" *)
  wire [15:0] REG_le_190;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:611" *)
  wire [15:0] REG_le_191;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:612" *)
  wire [15:0] REG_le_192;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:613" *)
  wire [15:0] REG_le_193;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:614" *)
  wire [15:0] REG_le_194;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:615" *)
  wire [15:0] REG_le_195;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:616" *)
  wire [15:0] REG_le_196;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:617" *)
  wire [15:0] REG_le_197;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:618" *)
  wire [15:0] REG_le_198;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:619" *)
  wire [15:0] REG_le_199;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:101" *)
  reg [15:0] REG_le_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:102" *)
  reg [15:0] REG_le_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:620" *)
  wire [15:0] REG_le_200;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:621" *)
  wire [15:0] REG_le_201;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:622" *)
  wire [15:0] REG_le_202;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:623" *)
  wire [15:0] REG_le_203;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:624" *)
  wire [15:0] REG_le_204;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:625" *)
  wire [15:0] REG_le_205;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:626" *)
  wire [15:0] REG_le_206;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:627" *)
  wire [15:0] REG_le_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:628" *)
  wire [15:0] REG_le_208;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:629" *)
  wire [15:0] REG_le_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:103" *)
  reg [15:0] REG_le_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:630" *)
  wire [15:0] REG_le_210;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:631" *)
  wire [15:0] REG_le_211;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:632" *)
  wire [15:0] REG_le_212;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:633" *)
  wire [15:0] REG_le_213;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:634" *)
  wire [15:0] REG_le_214;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:635" *)
  wire [15:0] REG_le_215;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:636" *)
  wire [15:0] REG_le_216;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:637" *)
  wire [15:0] REG_le_217;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:638" *)
  wire [15:0] REG_le_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:639" *)
  wire [15:0] REG_le_219;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:104" *)
  reg [15:0] REG_le_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:640" *)
  wire [15:0] REG_le_220;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:641" *)
  wire [15:0] REG_le_221;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:642" *)
  wire [15:0] REG_le_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:643" *)
  wire [15:0] REG_le_223;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:644" *)
  wire [15:0] REG_le_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:645" *)
  wire [15:0] REG_le_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:646" *)
  wire [15:0] REG_le_226;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:647" *)
  wire [15:0] REG_le_227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:648" *)
  wire [15:0] REG_le_228;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:649" *)
  wire [15:0] REG_le_229;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:105" *)
  reg [15:0] REG_le_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:650" *)
  wire [15:0] REG_le_230;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:651" *)
  wire [15:0] REG_le_231;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:652" *)
  wire [15:0] REG_le_232;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:653" *)
  wire [15:0] REG_le_233;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:654" *)
  wire [15:0] REG_le_234;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:655" *)
  wire [15:0] REG_le_235;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:656" *)
  wire [15:0] REG_le_236;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:657" *)
  wire [15:0] REG_le_237;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:658" *)
  wire [15:0] REG_le_238;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:659" *)
  wire [15:0] REG_le_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:106" *)
  reg [15:0] REG_le_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:660" *)
  wire [15:0] REG_le_240;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:661" *)
  wire [15:0] REG_le_241;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:662" *)
  wire [15:0] REG_le_242;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:663" *)
  wire [15:0] REG_le_243;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:664" *)
  wire [15:0] REG_le_244;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:665" *)
  wire [15:0] REG_le_245;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:666" *)
  wire [15:0] REG_le_246;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:667" *)
  wire [15:0] REG_le_247;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:668" *)
  wire [15:0] REG_le_248;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:669" *)
  wire [15:0] REG_le_249;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:107" *)
  reg [15:0] REG_le_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:670" *)
  wire [15:0] REG_le_250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:671" *)
  wire [15:0] REG_le_251;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:672" *)
  wire [15:0] REG_le_252;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:673" *)
  wire [15:0] REG_le_253;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:674" *)
  wire [15:0] REG_le_254;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:675" *)
  wire [15:0] REG_le_255;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:676" *)
  wire [15:0] REG_le_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:108" *)
  reg [15:0] REG_le_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:109" *)
  reg [15:0] REG_le_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:110" *)
  reg [15:0] REG_le_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:111" *)
  reg [15:0] REG_le_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:112" *)
  reg [15:0] REG_le_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:113" *)
  reg [15:0] REG_le_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:114" *)
  reg [15:0] REG_le_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:115" *)
  reg [15:0] REG_le_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:116" *)
  reg [15:0] REG_le_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:117" *)
  reg [15:0] REG_le_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:118" *)
  reg [15:0] REG_le_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:119" *)
  reg [15:0] REG_le_36;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:120" *)
  reg [15:0] REG_le_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:121" *)
  reg [15:0] REG_le_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:122" *)
  reg [15:0] REG_le_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:123" *)
  reg [15:0] REG_le_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:124" *)
  reg [15:0] REG_le_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:125" *)
  reg [15:0] REG_le_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:126" *)
  reg [15:0] REG_le_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:127" *)
  reg [15:0] REG_le_43;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:128" *)
  reg [15:0] REG_le_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:129" *)
  reg [15:0] REG_le_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:130" *)
  reg [15:0] REG_le_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:131" *)
  reg [15:0] REG_le_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:132" *)
  reg [15:0] REG_le_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:133" *)
  reg [15:0] REG_le_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:134" *)
  reg [15:0] REG_le_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:135" *)
  reg [15:0] REG_le_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:136" *)
  reg [15:0] REG_le_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:137" *)
  reg [15:0] REG_le_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:138" *)
  reg [15:0] REG_le_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:139" *)
  reg [15:0] REG_le_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:140" *)
  reg [15:0] REG_le_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:141" *)
  reg [15:0] REG_le_56;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:142" *)
  reg [15:0] REG_le_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:143" *)
  reg [15:0] REG_le_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:144" *)
  reg [15:0] REG_le_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:145" *)
  reg [15:0] REG_le_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:146" *)
  reg [15:0] REG_le_60;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:147" *)
  reg [15:0] REG_le_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:148" *)
  reg [15:0] REG_le_62;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:149" *)
  reg [15:0] REG_le_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:150" *)
  reg [15:0] REG_le_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:677" *)
  wire [15:0] REG_le_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:678" *)
  wire [15:0] REG_le_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:679" *)
  wire [15:0] REG_le_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:680" *)
  wire [15:0] REG_le_68;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:681" *)
  wire [15:0] REG_le_69;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:151" *)
  reg [15:0] REG_le_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:682" *)
  wire [15:0] REG_le_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:683" *)
  wire [15:0] REG_le_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:684" *)
  wire [15:0] REG_le_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:685" *)
  wire [15:0] REG_le_73;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:686" *)
  wire [15:0] REG_le_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:687" *)
  wire [15:0] REG_le_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:688" *)
  wire [15:0] REG_le_76;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:689" *)
  wire [15:0] REG_le_77;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:690" *)
  wire [15:0] REG_le_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:691" *)
  wire [15:0] REG_le_79;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:152" *)
  reg [15:0] REG_le_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:692" *)
  wire [15:0] REG_le_80;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:693" *)
  wire [15:0] REG_le_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:694" *)
  wire [15:0] REG_le_82;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:695" *)
  wire [15:0] REG_le_83;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:696" *)
  wire [15:0] REG_le_84;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:697" *)
  wire [15:0] REG_le_85;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:698" *)
  wire [15:0] REG_le_86;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:699" *)
  wire [15:0] REG_le_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:700" *)
  wire [15:0] REG_le_88;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:701" *)
  wire [15:0] REG_le_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:153" *)
  reg [15:0] REG_le_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:702" *)
  wire [15:0] REG_le_90;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:703" *)
  wire [15:0] REG_le_91;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:704" *)
  wire [15:0] REG_le_92;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:705" *)
  wire [15:0] REG_le_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:706" *)
  wire [15:0] REG_le_94;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:707" *)
  wire [15:0] REG_le_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:708" *)
  wire [15:0] REG_le_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:709" *)
  wire [15:0] REG_le_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:710" *)
  wire [15:0] REG_le_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:711" *)
  wire [15:0] REG_le_99;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:154" *)
  reg [15:0] REG_lo_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:155" *)
  reg [15:0] REG_lo_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:156" *)
  reg [15:0] REG_lo_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:157" *)
  reg [15:0] REG_lo_100;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:158" *)
  reg [15:0] REG_lo_101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:159" *)
  reg [15:0] REG_lo_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:160" *)
  reg [15:0] REG_lo_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:161" *)
  reg [15:0] REG_lo_104;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:162" *)
  reg [15:0] REG_lo_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:163" *)
  reg [15:0] REG_lo_106;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:164" *)
  reg [15:0] REG_lo_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:165" *)
  reg [15:0] REG_lo_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:166" *)
  reg [15:0] REG_lo_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:167" *)
  reg [15:0] REG_lo_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:168" *)
  reg [15:0] REG_lo_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:169" *)
  reg [15:0] REG_lo_111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:170" *)
  reg [15:0] REG_lo_112;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:171" *)
  reg [15:0] REG_lo_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:172" *)
  reg [15:0] REG_lo_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:173" *)
  reg [15:0] REG_lo_115;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:174" *)
  reg [15:0] REG_lo_116;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:175" *)
  reg [15:0] REG_lo_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:176" *)
  reg [15:0] REG_lo_118;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:177" *)
  reg [15:0] REG_lo_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:178" *)
  reg [15:0] REG_lo_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:179" *)
  reg [15:0] REG_lo_120;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:180" *)
  reg [15:0] REG_lo_121;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:181" *)
  reg [15:0] REG_lo_122;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:182" *)
  reg [15:0] REG_lo_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:183" *)
  reg [15:0] REG_lo_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:184" *)
  reg [15:0] REG_lo_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:185" *)
  reg [15:0] REG_lo_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:186" *)
  reg [15:0] REG_lo_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:187" *)
  reg [15:0] REG_lo_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:188" *)
  reg [15:0] REG_lo_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:189" *)
  reg [15:0] REG_lo_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:190" *)
  reg [15:0] REG_lo_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:191" *)
  reg [15:0] REG_lo_131;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:192" *)
  reg [15:0] REG_lo_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:193" *)
  reg [15:0] REG_lo_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:194" *)
  reg [15:0] REG_lo_134;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:195" *)
  reg [15:0] REG_lo_135;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:196" *)
  reg [15:0] REG_lo_136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:197" *)
  reg [15:0] REG_lo_137;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:198" *)
  reg [15:0] REG_lo_138;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:199" *)
  reg [15:0] REG_lo_139;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:200" *)
  reg [15:0] REG_lo_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:201" *)
  reg [15:0] REG_lo_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:202" *)
  reg [15:0] REG_lo_141;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:203" *)
  reg [15:0] REG_lo_142;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:204" *)
  reg [15:0] REG_lo_143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:205" *)
  reg [15:0] REG_lo_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:206" *)
  reg [15:0] REG_lo_145;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:207" *)
  reg [15:0] REG_lo_146;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:208" *)
  reg [15:0] REG_lo_147;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:209" *)
  reg [15:0] REG_lo_148;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:210" *)
  reg [15:0] REG_lo_149;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:211" *)
  reg [15:0] REG_lo_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:212" *)
  reg [15:0] REG_lo_150;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:213" *)
  reg [15:0] REG_lo_151;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:214" *)
  reg [15:0] REG_lo_152;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:215" *)
  reg [15:0] REG_lo_153;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:216" *)
  reg [15:0] REG_lo_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:217" *)
  reg [15:0] REG_lo_155;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:218" *)
  reg [15:0] REG_lo_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:219" *)
  reg [15:0] REG_lo_157;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:220" *)
  reg [15:0] REG_lo_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:221" *)
  reg [15:0] REG_lo_159;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:222" *)
  reg [15:0] REG_lo_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:223" *)
  reg [15:0] REG_lo_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:224" *)
  reg [15:0] REG_lo_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:225" *)
  reg [15:0] REG_lo_162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:226" *)
  reg [15:0] REG_lo_163;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:227" *)
  reg [15:0] REG_lo_164;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:228" *)
  reg [15:0] REG_lo_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:229" *)
  reg [15:0] REG_lo_166;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:230" *)
  reg [15:0] REG_lo_167;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:231" *)
  reg [15:0] REG_lo_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:232" *)
  reg [15:0] REG_lo_169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:233" *)
  reg [15:0] REG_lo_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:234" *)
  reg [15:0] REG_lo_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:235" *)
  reg [15:0] REG_lo_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:236" *)
  reg [15:0] REG_lo_172;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:237" *)
  reg [15:0] REG_lo_173;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:238" *)
  reg [15:0] REG_lo_174;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:239" *)
  reg [15:0] REG_lo_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:240" *)
  reg [15:0] REG_lo_176;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:241" *)
  reg [15:0] REG_lo_177;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:242" *)
  reg [15:0] REG_lo_178;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:243" *)
  reg [15:0] REG_lo_179;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:244" *)
  reg [15:0] REG_lo_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:245" *)
  reg [15:0] REG_lo_180;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:246" *)
  reg [15:0] REG_lo_181;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:247" *)
  reg [15:0] REG_lo_182;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:248" *)
  reg [15:0] REG_lo_183;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:249" *)
  reg [15:0] REG_lo_184;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:250" *)
  reg [15:0] REG_lo_185;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:251" *)
  reg [15:0] REG_lo_186;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:252" *)
  reg [15:0] REG_lo_187;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:253" *)
  reg [15:0] REG_lo_188;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:254" *)
  reg [15:0] REG_lo_189;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:255" *)
  reg [15:0] REG_lo_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:256" *)
  reg [15:0] REG_lo_190;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:257" *)
  reg [15:0] REG_lo_191;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:258" *)
  reg [15:0] REG_lo_192;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:259" *)
  reg [15:0] REG_lo_193;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:260" *)
  reg [15:0] REG_lo_194;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:261" *)
  reg [15:0] REG_lo_195;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:262" *)
  reg [15:0] REG_lo_196;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:263" *)
  reg [15:0] REG_lo_197;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:264" *)
  reg [15:0] REG_lo_198;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:265" *)
  reg [15:0] REG_lo_199;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:266" *)
  reg [15:0] REG_lo_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:267" *)
  reg [15:0] REG_lo_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:268" *)
  reg [15:0] REG_lo_200;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:269" *)
  reg [15:0] REG_lo_201;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:270" *)
  reg [15:0] REG_lo_202;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:271" *)
  reg [15:0] REG_lo_203;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:272" *)
  reg [15:0] REG_lo_204;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:273" *)
  reg [15:0] REG_lo_205;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:274" *)
  reg [15:0] REG_lo_206;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:275" *)
  reg [15:0] REG_lo_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:276" *)
  reg [15:0] REG_lo_208;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:277" *)
  reg [15:0] REG_lo_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:278" *)
  reg [15:0] REG_lo_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:279" *)
  reg [15:0] REG_lo_210;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:280" *)
  reg [15:0] REG_lo_211;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:281" *)
  reg [15:0] REG_lo_212;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:282" *)
  reg [15:0] REG_lo_213;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:283" *)
  reg [15:0] REG_lo_214;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:284" *)
  reg [15:0] REG_lo_215;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:285" *)
  reg [15:0] REG_lo_216;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:286" *)
  reg [15:0] REG_lo_217;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:287" *)
  reg [15:0] REG_lo_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:288" *)
  reg [15:0] REG_lo_219;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:289" *)
  reg [15:0] REG_lo_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:290" *)
  reg [15:0] REG_lo_220;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:291" *)
  reg [15:0] REG_lo_221;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:292" *)
  reg [15:0] REG_lo_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:293" *)
  reg [15:0] REG_lo_223;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:294" *)
  reg [15:0] REG_lo_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:295" *)
  reg [15:0] REG_lo_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:296" *)
  reg [15:0] REG_lo_226;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:297" *)
  reg [15:0] REG_lo_227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:298" *)
  reg [15:0] REG_lo_228;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:299" *)
  reg [15:0] REG_lo_229;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:300" *)
  reg [15:0] REG_lo_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:301" *)
  reg [15:0] REG_lo_230;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:302" *)
  reg [15:0] REG_lo_231;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:303" *)
  reg [15:0] REG_lo_232;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:304" *)
  reg [15:0] REG_lo_233;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:305" *)
  reg [15:0] REG_lo_234;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:306" *)
  reg [15:0] REG_lo_235;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:307" *)
  reg [15:0] REG_lo_236;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:308" *)
  reg [15:0] REG_lo_237;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:309" *)
  reg [15:0] REG_lo_238;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:310" *)
  reg [15:0] REG_lo_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:311" *)
  reg [15:0] REG_lo_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:312" *)
  reg [15:0] REG_lo_240;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:313" *)
  reg [15:0] REG_lo_241;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:314" *)
  reg [15:0] REG_lo_242;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:315" *)
  reg [15:0] REG_lo_243;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:316" *)
  reg [15:0] REG_lo_244;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:317" *)
  reg [15:0] REG_lo_245;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:318" *)
  reg [15:0] REG_lo_246;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:319" *)
  reg [15:0] REG_lo_247;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:320" *)
  reg [15:0] REG_lo_248;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:321" *)
  reg [15:0] REG_lo_249;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:322" *)
  reg [15:0] REG_lo_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:323" *)
  reg [15:0] REG_lo_250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:324" *)
  reg [15:0] REG_lo_251;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:325" *)
  reg [15:0] REG_lo_252;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:326" *)
  reg [15:0] REG_lo_253;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:327" *)
  reg [15:0] REG_lo_254;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:328" *)
  reg [15:0] REG_lo_255;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:329" *)
  reg [15:0] REG_lo_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:330" *)
  reg [15:0] REG_lo_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:331" *)
  reg [15:0] REG_lo_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:332" *)
  reg [15:0] REG_lo_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:333" *)
  reg [15:0] REG_lo_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:334" *)
  reg [15:0] REG_lo_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:335" *)
  reg [15:0] REG_lo_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:336" *)
  reg [15:0] REG_lo_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:337" *)
  reg [15:0] REG_lo_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:338" *)
  reg [15:0] REG_lo_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:339" *)
  reg [15:0] REG_lo_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:340" *)
  reg [15:0] REG_lo_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:341" *)
  reg [15:0] REG_lo_36;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:342" *)
  reg [15:0] REG_lo_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:343" *)
  reg [15:0] REG_lo_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:344" *)
  reg [15:0] REG_lo_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:345" *)
  reg [15:0] REG_lo_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:346" *)
  reg [15:0] REG_lo_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:347" *)
  reg [15:0] REG_lo_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:348" *)
  reg [15:0] REG_lo_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:349" *)
  reg [15:0] REG_lo_43;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:350" *)
  reg [15:0] REG_lo_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:351" *)
  reg [15:0] REG_lo_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:352" *)
  reg [15:0] REG_lo_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:353" *)
  reg [15:0] REG_lo_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:354" *)
  reg [15:0] REG_lo_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:355" *)
  reg [15:0] REG_lo_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:356" *)
  reg [15:0] REG_lo_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:357" *)
  reg [15:0] REG_lo_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:358" *)
  reg [15:0] REG_lo_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:359" *)
  reg [15:0] REG_lo_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:360" *)
  reg [15:0] REG_lo_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:361" *)
  reg [15:0] REG_lo_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:362" *)
  reg [15:0] REG_lo_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:363" *)
  reg [15:0] REG_lo_56;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:364" *)
  reg [15:0] REG_lo_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:365" *)
  reg [15:0] REG_lo_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:366" *)
  reg [15:0] REG_lo_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:367" *)
  reg [15:0] REG_lo_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:368" *)
  reg [15:0] REG_lo_60;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:369" *)
  reg [15:0] REG_lo_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:370" *)
  reg [15:0] REG_lo_62;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:371" *)
  reg [15:0] REG_lo_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:372" *)
  reg [15:0] REG_lo_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:373" *)
  reg [15:0] REG_lo_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:374" *)
  reg [15:0] REG_lo_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:375" *)
  reg [15:0] REG_lo_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:376" *)
  reg [15:0] REG_lo_68;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:377" *)
  reg [15:0] REG_lo_69;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:378" *)
  reg [15:0] REG_lo_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:379" *)
  reg [15:0] REG_lo_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:380" *)
  reg [15:0] REG_lo_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:381" *)
  reg [15:0] REG_lo_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:382" *)
  reg [15:0] REG_lo_73;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:383" *)
  reg [15:0] REG_lo_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:384" *)
  reg [15:0] REG_lo_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:385" *)
  reg [15:0] REG_lo_76;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:386" *)
  reg [15:0] REG_lo_77;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:387" *)
  reg [15:0] REG_lo_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:388" *)
  reg [15:0] REG_lo_79;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:389" *)
  reg [15:0] REG_lo_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:390" *)
  reg [15:0] REG_lo_80;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:391" *)
  reg [15:0] REG_lo_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:392" *)
  reg [15:0] REG_lo_82;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:393" *)
  reg [15:0] REG_lo_83;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:394" *)
  reg [15:0] REG_lo_84;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:395" *)
  reg [15:0] REG_lo_85;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:396" *)
  reg [15:0] REG_lo_86;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:397" *)
  reg [15:0] REG_lo_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:398" *)
  reg [15:0] REG_lo_88;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:399" *)
  reg [15:0] REG_lo_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:400" *)
  reg [15:0] REG_lo_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:401" *)
  reg [15:0] REG_lo_90;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:402" *)
  reg [15:0] REG_lo_91;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:403" *)
  reg [15:0] REG_lo_92;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:404" *)
  reg [15:0] REG_lo_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:405" *)
  reg [15:0] REG_lo_94;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:406" *)
  reg [15:0] REG_lo_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:407" *)
  reg [15:0] REG_lo_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:408" *)
  reg [15:0] REG_lo_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:409" *)
  reg [15:0] REG_lo_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:410" *)
  reg [15:0] REG_lo_99;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:712" *)
  wire [279:0] cmd_fifo_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:713" *)
  wire cmd_fifo_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:714" *)
  (* unused_bits = "0" *)
  wire cmd_fifo_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:715" *)
  wire [279:0] cmd_fifo_wr_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:716" *)
  wire cmd_fifo_wr_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:717" *)
  wire cmd_fifo_wr_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:718" *)
  wire [127:0] dat_fifo_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:719" *)
  wire dat_fifo_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:720" *)
  wire dat_fifo_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:721" *)
  wire [127:0] dat_fifo_wr_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:722" *)
  wire dat_fifo_wr_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:723" *)
  wire [15:0] dat_in_y0_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:724" *)
  wire [15:0] dat_in_y0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:725" *)
  wire [15:0] dat_in_y0_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:726" *)
  wire [15:0] dat_in_y0_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:727" *)
  wire [15:0] dat_in_y1_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:728" *)
  wire [15:0] dat_in_y1_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:729" *)
  wire [15:0] dat_in_y1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:730" *)
  wire [15:0] dat_in_y1_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:81" *)
  output [31:0] dp2reg_lut_hybrid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:82" *)
  output [15:0] dp2reg_lut_int_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:83" *)
  output [31:0] dp2reg_lut_le_hit;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:84" *)
  output [31:0] dp2reg_lut_lo_hit;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:85" *)
  output [31:0] dp2reg_lut_oflow;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:86" *)
  output [31:0] dp2reg_lut_uflow;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:59" *)
  input [323:0] idx2lut_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:58" *)
  output idx2lut_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:57" *)
  input idx2lut_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:412" *)
  wire [15:0] le_data0_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:413" *)
  wire [15:0] le_data0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:414" *)
  wire [15:0] le_data0_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:415" *)
  wire [15:0] le_data0_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:416" *)
  wire [15:0] le_data1_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:417" *)
  wire [15:0] le_data1_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:418" *)
  wire [15:0] le_data1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:419" *)
  wire [15:0] le_data1_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:420" *)
  wire [15:0] le_lut_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:731" *)
  wire le_wr_en_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:732" *)
  wire le_wr_en_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:733" *)
  wire le_wr_en_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:734" *)
  wire le_wr_en_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:735" *)
  wire le_wr_en_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:736" *)
  wire le_wr_en_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:737" *)
  wire le_wr_en_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:738" *)
  wire le_wr_en_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:739" *)
  wire le_wr_en_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:740" *)
  wire le_wr_en_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:741" *)
  wire le_wr_en_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:742" *)
  wire le_wr_en_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:743" *)
  wire le_wr_en_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:744" *)
  wire le_wr_en_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:745" *)
  wire le_wr_en_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:746" *)
  wire le_wr_en_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:747" *)
  wire le_wr_en_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:748" *)
  wire le_wr_en_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:749" *)
  wire le_wr_en_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:750" *)
  wire le_wr_en_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:751" *)
  wire le_wr_en_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:752" *)
  wire le_wr_en_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:753" *)
  wire le_wr_en_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:754" *)
  wire le_wr_en_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:755" *)
  wire le_wr_en_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:756" *)
  wire le_wr_en_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:757" *)
  wire le_wr_en_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:758" *)
  wire le_wr_en_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:759" *)
  wire le_wr_en_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:760" *)
  wire le_wr_en_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:761" *)
  wire le_wr_en_36;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:762" *)
  wire le_wr_en_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:763" *)
  wire le_wr_en_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:764" *)
  wire le_wr_en_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:765" *)
  wire le_wr_en_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:766" *)
  wire le_wr_en_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:767" *)
  wire le_wr_en_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:768" *)
  wire le_wr_en_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:769" *)
  wire le_wr_en_43;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:770" *)
  wire le_wr_en_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:771" *)
  wire le_wr_en_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:772" *)
  wire le_wr_en_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:773" *)
  wire le_wr_en_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:774" *)
  wire le_wr_en_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:775" *)
  wire le_wr_en_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:776" *)
  wire le_wr_en_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:777" *)
  wire le_wr_en_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:778" *)
  wire le_wr_en_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:779" *)
  wire le_wr_en_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:780" *)
  wire le_wr_en_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:781" *)
  wire le_wr_en_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:782" *)
  wire le_wr_en_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:783" *)
  wire le_wr_en_56;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:784" *)
  wire le_wr_en_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:785" *)
  wire le_wr_en_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:786" *)
  wire le_wr_en_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:787" *)
  wire le_wr_en_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:788" *)
  wire le_wr_en_60;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:789" *)
  wire le_wr_en_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:790" *)
  wire le_wr_en_62;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:791" *)
  wire le_wr_en_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:792" *)
  wire le_wr_en_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:793" *)
  wire le_wr_en_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:794" *)
  wire le_wr_en_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:795" *)
  wire le_wr_en_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:421" *)
  wire [15:0] lo_data0_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:422" *)
  wire [15:0] lo_data0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:423" *)
  wire [15:0] lo_data0_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:424" *)
  wire [15:0] lo_data0_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:425" *)
  wire [15:0] lo_data1_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:426" *)
  wire [15:0] lo_data1_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:427" *)
  wire [15:0] lo_data1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:428" *)
  wire [15:0] lo_data1_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:429" *)
  wire [15:0] lo_lut_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:796" *)
  wire lo_wr_en_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:797" *)
  wire lo_wr_en_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:798" *)
  wire lo_wr_en_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:799" *)
  wire lo_wr_en_100;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:800" *)
  wire lo_wr_en_101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:801" *)
  wire lo_wr_en_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:802" *)
  wire lo_wr_en_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:803" *)
  wire lo_wr_en_104;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:804" *)
  wire lo_wr_en_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:805" *)
  wire lo_wr_en_106;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:806" *)
  wire lo_wr_en_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:807" *)
  wire lo_wr_en_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:808" *)
  wire lo_wr_en_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:809" *)
  wire lo_wr_en_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:810" *)
  wire lo_wr_en_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:811" *)
  wire lo_wr_en_111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:812" *)
  wire lo_wr_en_112;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:813" *)
  wire lo_wr_en_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:814" *)
  wire lo_wr_en_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:815" *)
  wire lo_wr_en_115;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:816" *)
  wire lo_wr_en_116;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:817" *)
  wire lo_wr_en_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:818" *)
  wire lo_wr_en_118;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:819" *)
  wire lo_wr_en_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:820" *)
  wire lo_wr_en_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:821" *)
  wire lo_wr_en_120;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:822" *)
  wire lo_wr_en_121;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:823" *)
  wire lo_wr_en_122;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:824" *)
  wire lo_wr_en_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:825" *)
  wire lo_wr_en_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:826" *)
  wire lo_wr_en_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:827" *)
  wire lo_wr_en_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:828" *)
  wire lo_wr_en_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:829" *)
  wire lo_wr_en_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:830" *)
  wire lo_wr_en_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:831" *)
  wire lo_wr_en_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:832" *)
  wire lo_wr_en_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:833" *)
  wire lo_wr_en_131;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:834" *)
  wire lo_wr_en_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:835" *)
  wire lo_wr_en_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:836" *)
  wire lo_wr_en_134;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:837" *)
  wire lo_wr_en_135;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:838" *)
  wire lo_wr_en_136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:839" *)
  wire lo_wr_en_137;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:840" *)
  wire lo_wr_en_138;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:841" *)
  wire lo_wr_en_139;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:842" *)
  wire lo_wr_en_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:843" *)
  wire lo_wr_en_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:844" *)
  wire lo_wr_en_141;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:845" *)
  wire lo_wr_en_142;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:846" *)
  wire lo_wr_en_143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:847" *)
  wire lo_wr_en_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:848" *)
  wire lo_wr_en_145;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:849" *)
  wire lo_wr_en_146;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:850" *)
  wire lo_wr_en_147;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:851" *)
  wire lo_wr_en_148;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:852" *)
  wire lo_wr_en_149;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:853" *)
  wire lo_wr_en_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:854" *)
  wire lo_wr_en_150;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:855" *)
  wire lo_wr_en_151;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:856" *)
  wire lo_wr_en_152;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:857" *)
  wire lo_wr_en_153;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:858" *)
  wire lo_wr_en_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:859" *)
  wire lo_wr_en_155;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:860" *)
  wire lo_wr_en_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:861" *)
  wire lo_wr_en_157;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:862" *)
  wire lo_wr_en_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:863" *)
  wire lo_wr_en_159;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:864" *)
  wire lo_wr_en_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:865" *)
  wire lo_wr_en_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:866" *)
  wire lo_wr_en_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:867" *)
  wire lo_wr_en_162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:868" *)
  wire lo_wr_en_163;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:869" *)
  wire lo_wr_en_164;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:870" *)
  wire lo_wr_en_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:871" *)
  wire lo_wr_en_166;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:872" *)
  wire lo_wr_en_167;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:873" *)
  wire lo_wr_en_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:874" *)
  wire lo_wr_en_169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:875" *)
  wire lo_wr_en_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:876" *)
  wire lo_wr_en_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:877" *)
  wire lo_wr_en_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:878" *)
  wire lo_wr_en_172;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:879" *)
  wire lo_wr_en_173;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:880" *)
  wire lo_wr_en_174;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:881" *)
  wire lo_wr_en_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:882" *)
  wire lo_wr_en_176;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:883" *)
  wire lo_wr_en_177;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:884" *)
  wire lo_wr_en_178;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:885" *)
  wire lo_wr_en_179;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:886" *)
  wire lo_wr_en_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:887" *)
  wire lo_wr_en_180;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:888" *)
  wire lo_wr_en_181;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:889" *)
  wire lo_wr_en_182;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:890" *)
  wire lo_wr_en_183;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:891" *)
  wire lo_wr_en_184;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:892" *)
  wire lo_wr_en_185;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:893" *)
  wire lo_wr_en_186;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:894" *)
  wire lo_wr_en_187;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:895" *)
  wire lo_wr_en_188;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:896" *)
  wire lo_wr_en_189;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:897" *)
  wire lo_wr_en_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:898" *)
  wire lo_wr_en_190;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:899" *)
  wire lo_wr_en_191;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:900" *)
  wire lo_wr_en_192;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:901" *)
  wire lo_wr_en_193;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:902" *)
  wire lo_wr_en_194;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:903" *)
  wire lo_wr_en_195;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:904" *)
  wire lo_wr_en_196;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:905" *)
  wire lo_wr_en_197;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:906" *)
  wire lo_wr_en_198;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:907" *)
  wire lo_wr_en_199;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:908" *)
  wire lo_wr_en_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:909" *)
  wire lo_wr_en_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:910" *)
  wire lo_wr_en_200;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:911" *)
  wire lo_wr_en_201;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:912" *)
  wire lo_wr_en_202;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:913" *)
  wire lo_wr_en_203;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:914" *)
  wire lo_wr_en_204;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:915" *)
  wire lo_wr_en_205;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:916" *)
  wire lo_wr_en_206;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:917" *)
  wire lo_wr_en_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:918" *)
  wire lo_wr_en_208;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:919" *)
  wire lo_wr_en_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:920" *)
  wire lo_wr_en_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:921" *)
  wire lo_wr_en_210;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:922" *)
  wire lo_wr_en_211;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:923" *)
  wire lo_wr_en_212;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:924" *)
  wire lo_wr_en_213;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:925" *)
  wire lo_wr_en_214;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:926" *)
  wire lo_wr_en_215;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:927" *)
  wire lo_wr_en_216;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:928" *)
  wire lo_wr_en_217;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:929" *)
  wire lo_wr_en_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:930" *)
  wire lo_wr_en_219;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:931" *)
  wire lo_wr_en_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:932" *)
  wire lo_wr_en_220;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:933" *)
  wire lo_wr_en_221;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:934" *)
  wire lo_wr_en_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:935" *)
  wire lo_wr_en_223;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:936" *)
  wire lo_wr_en_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:937" *)
  wire lo_wr_en_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:938" *)
  wire lo_wr_en_226;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:939" *)
  wire lo_wr_en_227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:940" *)
  wire lo_wr_en_228;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:941" *)
  wire lo_wr_en_229;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:942" *)
  wire lo_wr_en_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:943" *)
  wire lo_wr_en_230;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:944" *)
  wire lo_wr_en_231;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:945" *)
  wire lo_wr_en_232;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:946" *)
  wire lo_wr_en_233;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:947" *)
  wire lo_wr_en_234;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:948" *)
  wire lo_wr_en_235;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:949" *)
  wire lo_wr_en_236;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:950" *)
  wire lo_wr_en_237;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:951" *)
  wire lo_wr_en_238;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:952" *)
  wire lo_wr_en_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:953" *)
  wire lo_wr_en_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:954" *)
  wire lo_wr_en_240;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:955" *)
  wire lo_wr_en_241;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:956" *)
  wire lo_wr_en_242;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:957" *)
  wire lo_wr_en_243;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:958" *)
  wire lo_wr_en_244;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:959" *)
  wire lo_wr_en_245;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:960" *)
  wire lo_wr_en_246;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:961" *)
  wire lo_wr_en_247;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:962" *)
  wire lo_wr_en_248;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:963" *)
  wire lo_wr_en_249;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:964" *)
  wire lo_wr_en_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:965" *)
  wire lo_wr_en_250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:966" *)
  wire lo_wr_en_251;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:967" *)
  wire lo_wr_en_252;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:968" *)
  wire lo_wr_en_253;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:969" *)
  wire lo_wr_en_254;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:970" *)
  wire lo_wr_en_255;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:971" *)
  wire lo_wr_en_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:972" *)
  wire lo_wr_en_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:973" *)
  wire lo_wr_en_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:974" *)
  wire lo_wr_en_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:975" *)
  wire lo_wr_en_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:976" *)
  wire lo_wr_en_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:977" *)
  wire lo_wr_en_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:978" *)
  wire lo_wr_en_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:979" *)
  wire lo_wr_en_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:980" *)
  wire lo_wr_en_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:981" *)
  wire lo_wr_en_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:982" *)
  wire lo_wr_en_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:983" *)
  wire lo_wr_en_36;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:984" *)
  wire lo_wr_en_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:985" *)
  wire lo_wr_en_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:986" *)
  wire lo_wr_en_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:987" *)
  wire lo_wr_en_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:988" *)
  wire lo_wr_en_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:989" *)
  wire lo_wr_en_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:990" *)
  wire lo_wr_en_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:991" *)
  wire lo_wr_en_43;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:992" *)
  wire lo_wr_en_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:993" *)
  wire lo_wr_en_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:994" *)
  wire lo_wr_en_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:995" *)
  wire lo_wr_en_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:996" *)
  wire lo_wr_en_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:997" *)
  wire lo_wr_en_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:998" *)
  wire lo_wr_en_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:999" *)
  wire lo_wr_en_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1000" *)
  wire lo_wr_en_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1001" *)
  wire lo_wr_en_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1002" *)
  wire lo_wr_en_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1003" *)
  wire lo_wr_en_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1004" *)
  wire lo_wr_en_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1005" *)
  wire lo_wr_en_56;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1006" *)
  wire lo_wr_en_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1007" *)
  wire lo_wr_en_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1008" *)
  wire lo_wr_en_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1009" *)
  wire lo_wr_en_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1010" *)
  wire lo_wr_en_60;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1011" *)
  wire lo_wr_en_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1012" *)
  wire lo_wr_en_62;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1013" *)
  wire lo_wr_en_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1014" *)
  wire lo_wr_en_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1015" *)
  wire lo_wr_en_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1016" *)
  wire lo_wr_en_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1017" *)
  wire lo_wr_en_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1018" *)
  wire lo_wr_en_68;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1019" *)
  wire lo_wr_en_69;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1020" *)
  wire lo_wr_en_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1021" *)
  wire lo_wr_en_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1022" *)
  wire lo_wr_en_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1023" *)
  wire lo_wr_en_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1024" *)
  wire lo_wr_en_73;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1025" *)
  wire lo_wr_en_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1026" *)
  wire lo_wr_en_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1027" *)
  wire lo_wr_en_76;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1028" *)
  wire lo_wr_en_77;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1029" *)
  wire lo_wr_en_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1030" *)
  wire lo_wr_en_79;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1031" *)
  wire lo_wr_en_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1032" *)
  wire lo_wr_en_80;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1033" *)
  wire lo_wr_en_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1034" *)
  wire lo_wr_en_82;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1035" *)
  wire lo_wr_en_83;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1036" *)
  wire lo_wr_en_84;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1037" *)
  wire lo_wr_en_85;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1038" *)
  wire lo_wr_en_86;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1039" *)
  wire lo_wr_en_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1040" *)
  wire lo_wr_en_88;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1041" *)
  wire lo_wr_en_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1042" *)
  wire lo_wr_en_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1043" *)
  wire lo_wr_en_90;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1044" *)
  wire lo_wr_en_91;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1045" *)
  wire lo_wr_en_92;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1046" *)
  wire lo_wr_en_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1047" *)
  wire lo_wr_en_94;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1048" *)
  wire lo_wr_en_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1049" *)
  wire lo_wr_en_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1050" *)
  wire lo_wr_en_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1051" *)
  wire lo_wr_en_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1052" *)
  wire lo_wr_en_99;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:56" *)
  output [739:0] lut2inp_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:55" *)
  input lut2inp_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:54" *)
  output lut2inp_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1053" *)
  wire lut_access_type;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1054" *)
  wire [9:0] lut_addr;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1055" *)
  wire [15:0] lut_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:432" *)
  wire [31:0] lut_hybrid_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1056" *)
  wire [2:0] lut_hybrid_sum;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1057" *)
  wire [8:0] lut_in_addr0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1058" *)
  wire [8:0] lut_in_addr0_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1059" *)
  wire [8:0] lut_in_addr0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1060" *)
  wire [8:0] lut_in_addr1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1061" *)
  wire [8:0] lut_in_addr1_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1062" *)
  wire [8:0] lut_in_addr1_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1063" *)
  wire [8:0] lut_in_addr2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1064" *)
  wire [8:0] lut_in_addr2_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1065" *)
  wire [8:0] lut_in_addr2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1066" *)
  wire [8:0] lut_in_addr3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1067" *)
  wire [8:0] lut_in_addr3_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1068" *)
  wire [8:0] lut_in_addr3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1069" *)
  wire [34:0] lut_in_fraction0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1070" *)
  wire [34:0] lut_in_fraction1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1071" *)
  wire [34:0] lut_in_fraction2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1072" *)
  wire [34:0] lut_in_fraction3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1073" *)
  wire lut_in_hybrid0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1074" *)
  wire lut_in_hybrid1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1075" *)
  wire lut_in_hybrid2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1076" *)
  wire lut_in_hybrid3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1077" *)
  wire lut_in_le_hit0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1078" *)
  wire lut_in_le_hit1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1079" *)
  wire lut_in_le_hit2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1080" *)
  wire lut_in_le_hit3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1081" *)
  wire lut_in_lo_hit0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1082" *)
  wire lut_in_lo_hit1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1083" *)
  wire lut_in_lo_hit2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1084" *)
  wire lut_in_lo_hit3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1085" *)
  wire lut_in_oflow0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1086" *)
  wire lut_in_oflow1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1087" *)
  wire lut_in_oflow2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1088" *)
  wire lut_in_oflow3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:433" *)
  wire [323:0] lut_in_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1089" *)
  wire lut_in_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:434" *)
  wire lut_in_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1090" *)
  wire lut_in_sel0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1091" *)
  wire lut_in_sel1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1092" *)
  wire lut_in_sel2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1093" *)
  wire lut_in_sel3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1094" *)
  wire lut_in_uflow0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1095" *)
  wire lut_in_uflow1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1096" *)
  wire lut_in_uflow2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1097" *)
  wire lut_in_uflow3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1098" *)
  wire [31:0] lut_in_x0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1099" *)
  wire [31:0] lut_in_x1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1100" *)
  wire [31:0] lut_in_x2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1101" *)
  wire [31:0] lut_in_x3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:435" *)
  wire [31:0] lut_le_hit_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1102" *)
  wire [2:0] lut_le_hit_sum;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:436" *)
  wire [31:0] lut_lo_hit_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1103" *)
  wire [2:0] lut_lo_hit_sum;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:437" *)
  wire [31:0] lut_oflow_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1104" *)
  wire [2:0] lut_oflow_sum;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1105" *)
  wire [739:0] lut_out_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:438" *)
  wire lut_out_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1106" *)
  wire lut_out_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1107" *)
  wire [27:0] lut_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1108" *)
  wire lut_table_id;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:439" *)
  wire [31:0] lut_uflow_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1109" *)
  wire [2:0] lut_uflow_sum;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1110" *)
  (* unused_bits = "0" *)
  wire mon_cmd_fifo_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:52" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:53" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:88" *)
  input op_en_load;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:440" *)
  wire [31:0] out_bias0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:444" *)
  wire [31:0] out_bias1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:448" *)
  wire [31:0] out_bias2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:452" *)
  wire [31:0] out_bias3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1111" *)
  wire out_flow0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1112" *)
  wire out_flow1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1113" *)
  wire out_flow2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1114" *)
  wire out_flow3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1115" *)
  wire [34:0] out_fraction0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1116" *)
  wire [34:0] out_fraction1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1117" *)
  wire [34:0] out_fraction2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1118" *)
  wire [34:0] out_fraction3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:456" *)
  wire [31:0] out_offset0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:457" *)
  wire [31:0] out_offset1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:458" *)
  wire [31:0] out_offset2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:459" *)
  wire [31:0] out_offset3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1119" *)
  wire out_oflow0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1120" *)
  wire out_oflow1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1121" *)
  wire out_oflow2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1122" *)
  wire out_oflow3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:460" *)
  wire [15:0] out_scale0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:461" *)
  wire [15:0] out_scale1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:462" *)
  wire [15:0] out_scale2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:463" *)
  wire [15:0] out_scale3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1123" *)
  wire out_sel0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1124" *)
  wire out_sel1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1125" *)
  wire out_sel2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1126" *)
  wire out_sel3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:464" *)
  wire [4:0] out_shift0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:465" *)
  wire [4:0] out_shift1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:466" *)
  wire [4:0] out_shift2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:467" *)
  wire [4:0] out_shift3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1127" *)
  wire out_uflow0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1128" *)
  wire out_uflow1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1129" *)
  wire out_uflow2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1130" *)
  wire out_uflow3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1131" *)
  wire [31:0] out_x0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1132" *)
  wire [31:0] out_x1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1133" *)
  wire [31:0] out_x2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1134" *)
  wire [31:0] out_x3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1135" *)
  wire [15:0] out_y0_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1136" *)
  wire [15:0] out_y0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1137" *)
  wire [15:0] out_y0_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1138" *)
  wire [15:0] out_y0_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1139" *)
  wire [15:0] out_y1_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1140" *)
  wire [15:0] out_y1_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1141" *)
  wire [15:0] out_y1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1142" *)
  wire [15:0] out_y1_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22250" *)
  wire p1_assert_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:468" *)
  reg [323:0] p1_pipe_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:469" *)
  wire [323:0] p1_pipe_rand_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:470" *)
  wire p1_pipe_rand_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:471" *)
  wire p1_pipe_rand_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:472" *)
  wire p1_pipe_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:473" *)
  wire p1_pipe_ready_bc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:474" *)
  reg p1_pipe_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31652" *)
  wire p2_assert_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:475" *)
  reg [739:0] p2_pipe_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:476" *)
  wire [739:0] p2_pipe_rand_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:477" *)
  wire p2_pipe_rand_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:478" *)
  wire p2_pipe_rand_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:479" *)
  reg p2_pipe_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:480" *)
  wire p2_pipe_ready_bc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:481" *)
  wire [739:0] p2_pipe_skid_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:482" *)
  wire p2_pipe_skid_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:483" *)
  wire p2_pipe_skid_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:484" *)
  reg p2_pipe_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:485" *)
  wire p2_skid_catch;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:486" *)
  reg [739:0] p2_skid_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:487" *)
  wire p2_skid_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:488" *)
  wire p2_skid_ready_flop;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:489" *)
  reg p2_skid_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1143" *)
  wire [2:0] perf_lut_hybrid_add;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:490" *)
  wire perf_lut_hybrid_adv;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:491" *)
  reg [31:0] perf_lut_hybrid_cnt_cur;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:492" *)
  wire [33:0] perf_lut_hybrid_cnt_ext;
  wire [31:0] perf_lut_hybrid_cnt_mod;
  wire [31:0] perf_lut_hybrid_cnt_new;
  wire [31:0] perf_lut_hybrid_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1144" *)
  wire perf_lut_hybrid_sub;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1145" *)
  wire [2:0] perf_lut_le_hit_add;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:496" *)
  wire perf_lut_le_hit_adv;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:497" *)
  reg [31:0] perf_lut_le_hit_cnt_cur;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:498" *)
  wire [33:0] perf_lut_le_hit_cnt_ext;
  wire [31:0] perf_lut_le_hit_cnt_mod;
  wire [31:0] perf_lut_le_hit_cnt_new;
  wire [31:0] perf_lut_le_hit_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1146" *)
  wire perf_lut_le_hit_sub;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1147" *)
  wire [2:0] perf_lut_lo_hit_add;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:502" *)
  wire perf_lut_lo_hit_adv;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:503" *)
  reg [31:0] perf_lut_lo_hit_cnt_cur;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:504" *)
  wire [33:0] perf_lut_lo_hit_cnt_ext;
  wire [31:0] perf_lut_lo_hit_cnt_mod;
  wire [31:0] perf_lut_lo_hit_cnt_new;
  wire [31:0] perf_lut_lo_hit_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1148" *)
  wire perf_lut_lo_hit_sub;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1149" *)
  wire [2:0] perf_lut_oflow_add;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:508" *)
  wire perf_lut_oflow_adv;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:509" *)
  reg [31:0] perf_lut_oflow_cnt_cur;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:510" *)
  wire [33:0] perf_lut_oflow_cnt_ext;
  wire [31:0] perf_lut_oflow_cnt_mod;
  wire [31:0] perf_lut_oflow_cnt_new;
  wire [31:0] perf_lut_oflow_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1150" *)
  wire perf_lut_oflow_sub;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1151" *)
  wire [2:0] perf_lut_uflow_add;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:514" *)
  wire perf_lut_uflow_adv;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:515" *)
  reg [31:0] perf_lut_uflow_cnt_cur;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:516" *)
  wire [33:0] perf_lut_uflow_cnt_ext;
  wire [31:0] perf_lut_uflow_cnt_mod;
  wire [31:0] perf_lut_uflow_cnt_new;
  wire [31:0] perf_lut_uflow_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1152" *)
  wire perf_lut_uflow_sub;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1153" *)
  wire [27:0] pro2lut_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1154" *)
  wire pro2lut_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1155" *)
  wire [9:0] pro_in_addr;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1156" *)
  wire [15:0] pro_in_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1157" *)
  wire pro_in_select_le;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1158" *)
  wire pro_in_select_lo;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1159" *)
  wire pro_in_table_id;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1160" *)
  wire pro_in_wr;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1161" *)
  wire pro_in_wr_en;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:87" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1162" *)
  wire rd_lut_en;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:60" *)
  input reg2dp_lut_int_access_type;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:61" *)
  input [9:0] reg2dp_lut_int_addr;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:62" *)
  input [15:0] reg2dp_lut_int_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:63" *)
  input reg2dp_lut_int_data_wr;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:64" *)
  input reg2dp_lut_int_table_id;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:65" *)
  input [31:0] reg2dp_lut_le_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:66" *)
  input reg2dp_lut_le_function;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:67" *)
  input [7:0] reg2dp_lut_le_index_offset;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:68" *)
  input [15:0] reg2dp_lut_le_slope_oflow_scale;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:69" *)
  input [4:0] reg2dp_lut_le_slope_oflow_shift;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:70" *)
  input [15:0] reg2dp_lut_le_slope_uflow_scale;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:71" *)
  input [4:0] reg2dp_lut_le_slope_uflow_shift;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:72" *)
  input [31:0] reg2dp_lut_le_start;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:73" *)
  input [31:0] reg2dp_lut_lo_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:74" *)
  input [15:0] reg2dp_lut_lo_slope_oflow_scale;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:75" *)
  input [4:0] reg2dp_lut_lo_slope_oflow_shift;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:76" *)
  input [15:0] reg2dp_lut_lo_slope_uflow_scale;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:77" *)
  input [4:0] reg2dp_lut_lo_slope_uflow_shift;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:78" *)
  input [31:0] reg2dp_lut_lo_start;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:79" *)
  input reg2dp_perf_lut_en;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:80" *)
  input [1:0] reg2dp_proc_precision;
  assign _0376_ = p1_pipe_data[271] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22380" *) p1_pipe_data[270];
  assign _0377_ = _0376_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22380" *) p1_pipe_data[269];
  assign lut_oflow_sum = _0377_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22380" *) p1_pipe_data[268];
  assign perf_lut_oflow_cnt_mod = perf_lut_oflow_cnt_cur + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22401" *) perf_lut_oflow_add;
  assign _0378_ = p1_pipe_data[275] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22423" *) p1_pipe_data[274];
  assign _0379_ = _0378_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22423" *) p1_pipe_data[273];
  assign lut_uflow_sum = _0379_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22423" *) p1_pipe_data[272];
  assign perf_lut_uflow_cnt_mod = perf_lut_uflow_cnt_cur + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22444" *) perf_lut_uflow_add;
  assign _0380_ = lut_in_hybrid3 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22470" *) lut_in_hybrid2;
  assign _0381_ = _0380_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22470" *) lut_in_hybrid1;
  assign lut_hybrid_sum = _0381_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22470" *) lut_in_hybrid0;
  assign perf_lut_hybrid_cnt_mod = perf_lut_hybrid_cnt_cur + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22491" *) perf_lut_hybrid_add;
  assign _0382_ = p1_pipe_data[319] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22513" *) p1_pipe_data[318];
  assign _0383_ = _0382_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22513" *) p1_pipe_data[317];
  assign lut_le_hit_sum = _0383_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22513" *) p1_pipe_data[316];
  assign perf_lut_le_hit_cnt_mod = perf_lut_le_hit_cnt_cur + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22534" *) perf_lut_le_hit_add;
  assign _0384_ = p1_pipe_data[323] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22556" *) p1_pipe_data[322];
  assign _0385_ = _0384_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22556" *) p1_pipe_data[321];
  assign lut_lo_hit_sum = _0385_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22556" *) p1_pipe_data[320];
  assign perf_lut_lo_hit_cnt_mod = perf_lut_lo_hit_cnt_cur + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22577" *) perf_lut_lo_hit_add;
  assign lut_in_addr0_1 = p1_pipe_data[288:280] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22604" *) 1'b1;
  assign lut_in_addr1_1 = p1_pipe_data[297:289] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22605" *) 1'b1;
  assign lut_in_addr2_1 = p1_pipe_data[306:298] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22606" *) 1'b1;
  assign lut_in_addr3_1 = p1_pipe_data[315:307] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22607" *) 1'b1;
  assign _0322_ = $signed(reg2dp_lut_le_index_offset) + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31129" *) $signed(8'b01111111);
  assign _0386_ = pro_in_wr_en & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10056" *) reg2dp_lut_int_table_id;
  assign lo_wr_en_64 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10056" *) _0388_;
  assign lo_wr_en_65 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10118" *) _0389_;
  assign lo_wr_en_66 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10180" *) _0390_;
  assign lo_wr_en_67 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10242" *) _0391_;
  assign lo_wr_en_68 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10304" *) _0392_;
  assign lo_wr_en_69 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10366" *) _0393_;
  assign lo_wr_en_70 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10428" *) _0394_;
  assign lo_wr_en_71 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10490" *) _0395_;
  assign lo_wr_en_72 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10552" *) _0396_;
  assign lo_wr_en_73 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10614" *) _0397_;
  assign lo_wr_en_74 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10676" *) _0398_;
  assign lo_wr_en_75 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10738" *) _0399_;
  assign lo_wr_en_76 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10800" *) _0400_;
  assign lo_wr_en_77 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10862" *) _0401_;
  assign lo_wr_en_78 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10924" *) _0402_;
  assign lo_wr_en_79 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10986" *) _0403_;
  assign lo_wr_en_80 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11048" *) _0404_;
  assign lo_wr_en_81 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11110" *) _0405_;
  assign lo_wr_en_82 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11172" *) _0406_;
  assign lo_wr_en_83 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11234" *) _0407_;
  assign lo_wr_en_84 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11296" *) _0408_;
  assign lo_wr_en_85 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11358" *) _0409_;
  assign lo_wr_en_86 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11420" *) _0410_;
  assign lo_wr_en_87 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11482" *) _0411_;
  assign lo_wr_en_88 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11544" *) _0412_;
  assign lo_wr_en_89 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11606" *) _0413_;
  assign lo_wr_en_90 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11668" *) _0414_;
  assign lo_wr_en_91 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11730" *) _0415_;
  assign lo_wr_en_92 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11792" *) _0416_;
  assign lo_wr_en_93 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11854" *) _0417_;
  assign pro_in_wr_en = reg2dp_lut_int_data_wr & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1191" *) reg2dp_lut_int_access_type;
  assign lo_wr_en_94 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11916" *) _0418_;
  assign lo_wr_en_95 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11978" *) _0419_;
  assign lo_wr_en_96 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12040" *) _0420_;
  assign lo_wr_en_97 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12102" *) _0421_;
  assign lo_wr_en_98 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12164" *) _0422_;
  assign lo_wr_en_99 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12226" *) _0423_;
  assign lo_wr_en_100 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12288" *) _0424_;
  assign lo_wr_en_101 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12350" *) _0425_;
  assign lo_wr_en_102 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12412" *) _0426_;
  assign lo_wr_en_103 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12474" *) _0427_;
  assign lo_wr_en_104 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12536" *) _0428_;
  assign lo_wr_en_105 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12598" *) _0429_;
  assign lo_wr_en_106 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12660" *) _0430_;
  assign lo_wr_en_107 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12722" *) _0431_;
  assign lo_wr_en_108 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12784" *) _0432_;
  assign lo_wr_en_109 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12846" *) _0433_;
  assign lo_wr_en_110 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12908" *) _0434_;
  assign lo_wr_en_111 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12970" *) _0435_;
  assign lo_wr_en_112 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13032" *) _0436_;
  assign lo_wr_en_113 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13094" *) _0437_;
  assign lo_wr_en_114 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13156" *) _0438_;
  assign lo_wr_en_115 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13218" *) _0439_;
  assign lo_wr_en_116 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13280" *) _0440_;
  assign lo_wr_en_117 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13342" *) _0441_;
  assign lo_wr_en_118 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13404" *) _0442_;
  assign lo_wr_en_119 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13466" *) _0443_;
  assign lo_wr_en_120 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13528" *) _0444_;
  assign lo_wr_en_121 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13590" *) _0445_;
  assign lo_wr_en_122 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13652" *) _0446_;
  assign lo_wr_en_123 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13714" *) _0447_;
  assign lo_wr_en_124 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13776" *) _0448_;
  assign lo_wr_en_125 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13838" *) _0449_;
  assign lo_wr_en_126 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13900" *) _0450_;
  assign lo_wr_en_127 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13962" *) _0451_;
  assign lo_wr_en_128 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14024" *) _0452_;
  assign lo_wr_en_129 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14086" *) _0453_;
  assign lo_wr_en_130 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14148" *) _0454_;
  assign lo_wr_en_131 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14210" *) _0455_;
  assign lo_wr_en_132 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14272" *) _0456_;
  assign lo_wr_en_133 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14334" *) _0457_;
  assign lo_wr_en_134 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14396" *) _0458_;
  assign lo_wr_en_135 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14458" *) _0459_;
  assign lo_wr_en_136 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14520" *) _0460_;
  assign lo_wr_en_137 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14582" *) _0461_;
  assign lo_wr_en_138 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14644" *) _0462_;
  assign lo_wr_en_139 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14706" *) _0463_;
  assign lo_wr_en_140 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14768" *) _0464_;
  assign lo_wr_en_141 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14830" *) _0465_;
  assign lo_wr_en_142 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14892" *) _0466_;
  assign lo_wr_en_143 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14954" *) _0467_;
  assign lo_wr_en_144 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15016" *) _0468_;
  assign lo_wr_en_145 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15078" *) _0469_;
  assign lo_wr_en_146 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15140" *) _0470_;
  assign lo_wr_en_147 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15202" *) _0471_;
  assign lo_wr_en_148 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15264" *) _0472_;
  assign lo_wr_en_149 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15326" *) _0473_;
  assign lo_wr_en_150 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15388" *) _0474_;
  assign lo_wr_en_151 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15450" *) _0475_;
  assign lo_wr_en_152 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15512" *) _0476_;
  assign lo_wr_en_153 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15574" *) _0477_;
  assign lo_wr_en_154 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15636" *) _0478_;
  assign lo_wr_en_155 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15698" *) _0479_;
  assign lo_wr_en_156 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15760" *) _0480_;
  assign lo_wr_en_157 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15822" *) _0481_;
  assign lo_wr_en_158 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15884" *) _0482_;
  assign lo_wr_en_159 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15946" *) _0483_;
  assign lo_wr_en_160 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16008" *) _0484_;
  assign lo_wr_en_161 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16070" *) _0485_;
  assign lo_wr_en_162 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16132" *) _0486_;
  assign lo_wr_en_163 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16194" *) _0487_;
  assign lo_wr_en_164 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16256" *) _0488_;
  assign lo_wr_en_165 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16318" *) _0489_;
  assign lo_wr_en_166 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16380" *) _0490_;
  assign lo_wr_en_167 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16442" *) _0491_;
  assign lo_wr_en_168 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16504" *) _0492_;
  assign lo_wr_en_169 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16566" *) _0493_;
  assign lo_wr_en_170 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16628" *) _0494_;
  assign lo_wr_en_171 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16690" *) _0495_;
  assign lo_wr_en_172 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16752" *) _0496_;
  assign lo_wr_en_173 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16814" *) _0497_;
  assign lo_wr_en_174 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16876" *) _0498_;
  assign lo_wr_en_175 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16938" *) _0499_;
  assign lo_wr_en_176 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17000" *) _0500_;
  assign lo_wr_en_177 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17062" *) _0501_;
  assign lo_wr_en_178 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17124" *) _0502_;
  assign lo_wr_en_179 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17186" *) _0503_;
  assign lo_wr_en_180 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17248" *) _0504_;
  assign lo_wr_en_181 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17310" *) _0505_;
  assign lo_wr_en_182 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17372" *) _0506_;
  assign lo_wr_en_183 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17434" *) _0507_;
  assign lo_wr_en_184 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17496" *) _0508_;
  assign lo_wr_en_185 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17558" *) _0509_;
  assign lo_wr_en_186 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17620" *) _0510_;
  assign lo_wr_en_187 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17682" *) _0511_;
  assign lo_wr_en_188 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17744" *) _0512_;
  assign lo_wr_en_189 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17806" *) _0513_;
  assign lo_wr_en_190 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17868" *) _0514_;
  assign lo_wr_en_191 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17930" *) _0515_;
  assign lo_wr_en_192 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17992" *) _0516_;
  assign lo_wr_en_193 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18054" *) _0517_;
  assign lo_wr_en_194 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18116" *) _0518_;
  assign lo_wr_en_195 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18178" *) _0519_;
  assign lo_wr_en_196 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18240" *) _0520_;
  assign lo_wr_en_197 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18302" *) _0521_;
  assign lo_wr_en_198 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18364" *) _0522_;
  assign lo_wr_en_199 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18426" *) _0523_;
  assign lo_wr_en_200 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18488" *) _0524_;
  assign lo_wr_en_201 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18550" *) _0525_;
  assign lo_wr_en_202 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18612" *) _0526_;
  assign _0387_ = pro_in_wr_en & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1866" *) pro_in_select_le;
  assign le_wr_en_0 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1866" *) _0527_;
  assign lo_wr_en_203 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18674" *) _0528_;
  assign lo_wr_en_204 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18736" *) _0529_;
  assign lo_wr_en_205 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18798" *) _0530_;
  assign lo_wr_en_206 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18860" *) _0531_;
  assign lo_wr_en_207 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18922" *) _0532_;
  assign lo_wr_en_208 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18984" *) _0533_;
  assign lo_wr_en_209 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19046" *) _0534_;
  assign lo_wr_en_210 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19108" *) _0535_;
  assign lo_wr_en_211 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19170" *) _0536_;
  assign lo_wr_en_212 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19232" *) _0537_;
  assign le_wr_en_1 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1928" *) _0538_;
  assign lo_wr_en_213 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19294" *) _0539_;
  assign lo_wr_en_214 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19356" *) _0540_;
  assign lo_wr_en_215 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19418" *) _0541_;
  assign lo_wr_en_216 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19480" *) _0542_;
  assign lo_wr_en_217 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19542" *) _0543_;
  assign lo_wr_en_218 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19604" *) _0544_;
  assign lo_wr_en_219 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19666" *) _0545_;
  assign lo_wr_en_220 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19728" *) _0546_;
  assign lo_wr_en_221 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19790" *) _0547_;
  assign lo_wr_en_222 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19852" *) _0548_;
  assign le_wr_en_2 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1990" *) _0549_;
  assign lo_wr_en_223 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19914" *) _0550_;
  assign lo_wr_en_224 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19976" *) _0551_;
  assign lo_wr_en_225 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20038" *) _0552_;
  assign lo_wr_en_226 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20100" *) _0553_;
  assign lo_wr_en_227 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20162" *) _0554_;
  assign lo_wr_en_228 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20224" *) _0555_;
  assign lo_wr_en_229 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20286" *) _0556_;
  assign lo_wr_en_230 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20348" *) _0557_;
  assign lo_wr_en_231 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20410" *) _0558_;
  assign lo_wr_en_232 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20472" *) _0559_;
  assign le_wr_en_3 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2052" *) _0560_;
  assign lo_wr_en_233 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20534" *) _0561_;
  assign lo_wr_en_234 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20596" *) _0562_;
  assign lo_wr_en_235 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20658" *) _0563_;
  assign lo_wr_en_236 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20720" *) _0564_;
  assign lo_wr_en_237 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20782" *) _0565_;
  assign lo_wr_en_238 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20844" *) _0566_;
  assign lo_wr_en_239 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20906" *) _0567_;
  assign lo_wr_en_240 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20968" *) _0568_;
  assign lo_wr_en_241 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21030" *) _0569_;
  assign lo_wr_en_242 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21092" *) _0570_;
  assign le_wr_en_4 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2114" *) _0571_;
  assign lo_wr_en_243 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21154" *) _0572_;
  assign lo_wr_en_244 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21216" *) _0573_;
  assign lo_wr_en_245 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21278" *) _0574_;
  assign lo_wr_en_246 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21340" *) _0575_;
  assign lo_wr_en_247 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21402" *) _0576_;
  assign lo_wr_en_248 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21464" *) _0577_;
  assign lo_wr_en_249 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21526" *) _0578_;
  assign lo_wr_en_250 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21588" *) _0579_;
  assign lo_wr_en_251 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21650" *) _0580_;
  assign lo_wr_en_252 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21712" *) _0581_;
  assign le_wr_en_5 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2176" *) _0582_;
  assign lo_wr_en_253 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21774" *) _0583_;
  assign lo_wr_en_254 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21836" *) _0584_;
  assign lo_wr_en_255 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21898" *) _0585_;
  assign lo_wr_en_256 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21960" *) _0586_;
  assign le_wr_en_6 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2238" *) _0587_;
  assign le_wr_en_7 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2300" *) _0588_;
  assign le_wr_en_8 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2362" *) _0589_;
  assign le_wr_en_9 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2424" *) _0590_;
  assign le_wr_en_10 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2486" *) _0591_;
  assign le_wr_en_11 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2548" *) _0592_;
  assign le_wr_en_12 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2610" *) _0593_;
  assign le_wr_en_13 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2672" *) _0594_;
  assign le_wr_en_14 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2734" *) _0595_;
  assign le_wr_en_15 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2796" *) _0596_;
  assign le_wr_en_16 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2858" *) _0597_;
  assign le_wr_en_17 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2920" *) _0598_;
  assign le_wr_en_18 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2982" *) _0599_;
  assign le_wr_en_19 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3044" *) _0600_;
  assign dat_fifo_wr_pvld = p1_pipe_valid & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31002" *) cmd_fifo_wr_prdy;
  assign le_wr_en_20 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3106" *) _0601_;
  assign cmd_fifo_rd_prdy = dat_fifo_rd_prdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31063" *) dat_fifo_rd_pvld;
  assign le_wr_en_21 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3168" *) _0603_;
  assign le_wr_en_22 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3230" *) _0604_;
  assign le_wr_en_23 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3292" *) _0605_;
  assign le_wr_en_24 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3354" *) _0606_;
  assign le_wr_en_25 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3416" *) _0607_;
  assign le_wr_en_26 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3478" *) _0608_;
  assign le_wr_en_27 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3540" *) _0609_;
  assign le_wr_en_28 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3602" *) _0610_;
  assign le_wr_en_29 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3664" *) _0611_;
  assign le_wr_en_30 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3726" *) _0612_;
  assign le_wr_en_31 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3788" *) _0613_;
  assign le_wr_en_32 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3850" *) _0614_;
  assign le_wr_en_33 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3912" *) _0615_;
  assign le_wr_en_34 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3974" *) _0616_;
  assign le_wr_en_35 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4036" *) _0617_;
  assign le_wr_en_36 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4098" *) _0618_;
  assign le_wr_en_37 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4160" *) _0619_;
  assign le_wr_en_38 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4222" *) _0620_;
  assign le_wr_en_39 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4284" *) _0621_;
  assign le_wr_en_40 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4346" *) _0622_;
  assign le_wr_en_41 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4408" *) _0623_;
  assign le_wr_en_42 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4470" *) _0624_;
  assign le_wr_en_43 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4532" *) _0625_;
  assign le_wr_en_44 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4594" *) _0626_;
  assign le_wr_en_45 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4656" *) _0627_;
  assign le_wr_en_46 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4718" *) _0628_;
  assign le_wr_en_47 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4780" *) _0629_;
  assign le_wr_en_48 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4842" *) _0630_;
  assign le_wr_en_49 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4904" *) _0631_;
  assign le_wr_en_50 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4966" *) _0632_;
  assign le_wr_en_51 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5028" *) _0633_;
  assign le_wr_en_52 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5090" *) _0634_;
  assign le_wr_en_53 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5152" *) _0635_;
  assign le_wr_en_54 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5214" *) _0636_;
  assign le_wr_en_55 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5276" *) _0637_;
  assign le_wr_en_56 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5338" *) _0638_;
  assign le_wr_en_57 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5400" *) _0639_;
  assign le_wr_en_58 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5462" *) _0640_;
  assign le_wr_en_59 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5524" *) _0641_;
  assign le_wr_en_60 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5586" *) _0642_;
  assign le_wr_en_61 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5648" *) _0643_;
  assign le_wr_en_62 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5710" *) _0644_;
  assign le_wr_en_63 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5772" *) _0645_;
  assign le_wr_en_64 = _0387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5834" *) _0388_;
  assign lo_wr_en_0 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6088" *) _0527_;
  assign lo_wr_en_1 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6150" *) _0538_;
  assign lo_wr_en_2 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6212" *) _0549_;
  assign lo_wr_en_3 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6274" *) _0560_;
  assign lo_wr_en_4 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6336" *) _0571_;
  assign lo_wr_en_5 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6398" *) _0582_;
  assign lo_wr_en_6 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6460" *) _0587_;
  assign lo_wr_en_7 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6522" *) _0588_;
  assign lo_wr_en_8 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6584" *) _0589_;
  assign lo_wr_en_9 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6646" *) _0590_;
  assign lo_wr_en_10 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6708" *) _0591_;
  assign lo_wr_en_11 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6770" *) _0592_;
  assign lo_wr_en_12 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6832" *) _0593_;
  assign lo_wr_en_13 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6894" *) _0594_;
  assign lo_wr_en_14 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6956" *) _0595_;
  assign lo_wr_en_15 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7018" *) _0596_;
  assign lo_wr_en_16 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7080" *) _0597_;
  assign lo_wr_en_17 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7142" *) _0598_;
  assign lo_wr_en_18 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7204" *) _0599_;
  assign lo_wr_en_19 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7266" *) _0600_;
  assign lo_wr_en_20 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7328" *) _0601_;
  assign lo_wr_en_21 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7390" *) _0603_;
  assign lo_wr_en_22 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7452" *) _0604_;
  assign lo_wr_en_23 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7514" *) _0605_;
  assign lo_wr_en_24 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7576" *) _0606_;
  assign lo_wr_en_25 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7638" *) _0607_;
  assign lo_wr_en_26 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7700" *) _0608_;
  assign lo_wr_en_27 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7762" *) _0609_;
  assign lo_wr_en_28 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7824" *) _0610_;
  assign lo_wr_en_29 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7886" *) _0611_;
  assign lo_wr_en_30 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7948" *) _0612_;
  assign lo_wr_en_31 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8010" *) _0613_;
  assign lo_wr_en_32 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8072" *) _0614_;
  assign lo_wr_en_33 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8134" *) _0615_;
  assign lo_wr_en_34 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8196" *) _0616_;
  assign lo_wr_en_35 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8258" *) _0617_;
  assign lo_wr_en_36 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8320" *) _0618_;
  assign lo_wr_en_37 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8382" *) _0619_;
  assign lo_wr_en_38 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8444" *) _0620_;
  assign lo_wr_en_39 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8506" *) _0621_;
  assign lo_wr_en_40 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8568" *) _0622_;
  assign lo_wr_en_41 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8630" *) _0623_;
  assign lo_wr_en_42 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8692" *) _0624_;
  assign lo_wr_en_43 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8754" *) _0625_;
  assign lo_wr_en_44 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8816" *) _0626_;
  assign lo_wr_en_45 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8878" *) _0627_;
  assign lo_wr_en_46 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8940" *) _0628_;
  assign lo_wr_en_47 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9002" *) _0629_;
  assign lo_wr_en_48 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9064" *) _0630_;
  assign lo_wr_en_49 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9126" *) _0631_;
  assign lo_wr_en_50 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9188" *) _0632_;
  assign lo_wr_en_51 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9250" *) _0633_;
  assign lo_wr_en_52 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9312" *) _0634_;
  assign lo_wr_en_53 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9374" *) _0635_;
  assign lo_wr_en_54 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9436" *) _0636_;
  assign lo_wr_en_55 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9498" *) _0637_;
  assign lo_wr_en_56 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9560" *) _0638_;
  assign lo_wr_en_57 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9622" *) _0639_;
  assign lo_wr_en_58 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9684" *) _0640_;
  assign lo_wr_en_59 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9746" *) _0641_;
  assign lo_wr_en_60 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9808" *) _0642_;
  assign lo_wr_en_61 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9870" *) _0643_;
  assign lo_wr_en_62 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9932" *) _0644_;
  assign lo_wr_en_63 = _0386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9994" *) _0645_;
  assign _0388_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10056" *) 7'b1000000;
  assign _0389_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10118" *) 7'b1000001;
  assign _0390_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10180" *) 7'b1000010;
  assign _0391_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10242" *) 7'b1000011;
  assign _0392_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10304" *) 7'b1000100;
  assign _0393_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10366" *) 7'b1000101;
  assign _0394_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10428" *) 7'b1000110;
  assign _0395_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10490" *) 7'b1000111;
  assign _0396_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10552" *) 7'b1001000;
  assign _0397_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10614" *) 7'b1001001;
  assign _0398_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10676" *) 7'b1001010;
  assign _0399_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10738" *) 7'b1001011;
  assign _0400_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10800" *) 7'b1001100;
  assign _0401_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10862" *) 7'b1001101;
  assign _0402_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10924" *) 7'b1001110;
  assign _0403_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10986" *) 7'b1001111;
  assign _0404_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11048" *) 7'b1010000;
  assign _0405_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11110" *) 7'b1010001;
  assign _0406_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11172" *) 7'b1010010;
  assign _0407_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11234" *) 7'b1010011;
  assign _0408_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11296" *) 7'b1010100;
  assign _0409_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11358" *) 7'b1010101;
  assign _0410_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11420" *) 7'b1010110;
  assign _0411_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11482" *) 7'b1010111;
  assign _0412_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11544" *) 7'b1011000;
  assign _0413_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11606" *) 7'b1011001;
  assign _0414_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11668" *) 7'b1011010;
  assign _0415_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11730" *) 7'b1011011;
  assign _0416_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11792" *) 7'b1011100;
  assign _0417_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11854" *) 7'b1011101;
  assign _0418_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11916" *) 7'b1011110;
  assign pro_in_select_le = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1193" *) reg2dp_lut_int_table_id;
  assign _0419_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11978" *) 7'b1011111;
  assign _0420_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12040" *) 7'b1100000;
  assign _0421_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12102" *) 7'b1100001;
  assign _0422_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12164" *) 7'b1100010;
  assign _0423_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12226" *) 7'b1100011;
  assign _0424_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12288" *) 7'b1100100;
  assign _0425_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12350" *) 7'b1100101;
  assign _0426_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12412" *) 7'b1100110;
  assign _0427_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12474" *) 7'b1100111;
  assign _0428_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12536" *) 7'b1101000;
  assign _0429_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12598" *) 7'b1101001;
  assign _0430_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12660" *) 7'b1101010;
  assign _0431_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12722" *) 7'b1101011;
  assign _0432_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12784" *) 7'b1101100;
  assign _0433_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12846" *) 7'b1101101;
  assign _0434_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12908" *) 7'b1101110;
  assign _0435_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12970" *) 7'b1101111;
  assign _0436_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13032" *) 7'b1110000;
  assign _0437_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13094" *) 7'b1110001;
  assign _0438_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13156" *) 7'b1110010;
  assign _0439_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13218" *) 7'b1110011;
  assign _0440_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13280" *) 7'b1110100;
  assign _0441_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13342" *) 7'b1110101;
  assign _0442_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13404" *) 7'b1110110;
  assign _0443_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13466" *) 7'b1110111;
  assign _0444_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13528" *) 7'b1111000;
  assign _0445_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13590" *) 7'b1111001;
  assign _0446_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13652" *) 7'b1111010;
  assign _0447_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13714" *) 7'b1111011;
  assign _0448_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13776" *) 7'b1111100;
  assign _0449_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13838" *) 7'b1111101;
  assign _0450_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13900" *) 7'b1111110;
  assign _0451_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13962" *) 7'b1111111;
  assign _0452_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14024" *) 8'b10000000;
  assign _0453_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14086" *) 8'b10000001;
  assign _0454_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14148" *) 8'b10000010;
  assign _0455_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14210" *) 8'b10000011;
  assign _0456_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14272" *) 8'b10000100;
  assign _0457_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14334" *) 8'b10000101;
  assign _0458_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14396" *) 8'b10000110;
  assign _0459_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14458" *) 8'b10000111;
  assign _0460_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14520" *) 8'b10001000;
  assign _0461_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14582" *) 8'b10001001;
  assign _0462_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14644" *) 8'b10001010;
  assign _0463_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14706" *) 8'b10001011;
  assign _0464_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14768" *) 8'b10001100;
  assign _0465_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14830" *) 8'b10001101;
  assign _0466_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14892" *) 8'b10001110;
  assign _0467_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14954" *) 8'b10001111;
  assign _0468_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15016" *) 8'b10010000;
  assign _0469_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15078" *) 8'b10010001;
  assign _0470_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15140" *) 8'b10010010;
  assign _0471_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15202" *) 8'b10010011;
  assign _0472_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15264" *) 8'b10010100;
  assign _0473_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15326" *) 8'b10010101;
  assign _0474_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15388" *) 8'b10010110;
  assign _0475_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15450" *) 8'b10010111;
  assign _0476_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15512" *) 8'b10011000;
  assign _0477_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15574" *) 8'b10011001;
  assign _0478_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15636" *) 8'b10011010;
  assign _0479_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15698" *) 8'b10011011;
  assign _0480_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15760" *) 8'b10011100;
  assign _0481_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15822" *) 8'b10011101;
  assign _0482_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15884" *) 8'b10011110;
  assign _0483_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15946" *) 8'b10011111;
  assign _0484_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16008" *) 8'b10100000;
  assign _0485_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16070" *) 8'b10100001;
  assign _0486_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16132" *) 8'b10100010;
  assign _0487_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16194" *) 8'b10100011;
  assign _0488_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16256" *) 8'b10100100;
  assign _0489_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16318" *) 8'b10100101;
  assign _0490_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16380" *) 8'b10100110;
  assign _0491_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16442" *) 8'b10100111;
  assign _0492_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16504" *) 8'b10101000;
  assign _0493_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16566" *) 8'b10101001;
  assign _0494_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16628" *) 8'b10101010;
  assign _0495_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16690" *) 8'b10101011;
  assign _0496_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16752" *) 8'b10101100;
  assign _0497_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16814" *) 8'b10101101;
  assign _0498_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16876" *) 8'b10101110;
  assign _0499_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16938" *) 8'b10101111;
  assign _0500_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17000" *) 8'b10110000;
  assign _0501_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17062" *) 8'b10110001;
  assign _0502_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17124" *) 8'b10110010;
  assign _0503_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17186" *) 8'b10110011;
  assign _0504_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17248" *) 8'b10110100;
  assign _0505_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17310" *) 8'b10110101;
  assign _0506_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17372" *) 8'b10110110;
  assign _0507_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17434" *) 8'b10110111;
  assign _0508_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17496" *) 8'b10111000;
  assign _0509_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17558" *) 8'b10111001;
  assign _0510_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17620" *) 8'b10111010;
  assign _0511_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17682" *) 8'b10111011;
  assign _0512_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17744" *) 8'b10111100;
  assign _0513_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17806" *) 8'b10111101;
  assign _0514_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17868" *) 8'b10111110;
  assign _0515_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17930" *) 8'b10111111;
  assign _0516_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17992" *) 8'b11000000;
  assign _0517_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18054" *) 8'b11000001;
  assign _0518_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18116" *) 8'b11000010;
  assign _0519_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18178" *) 8'b11000011;
  assign _0520_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18240" *) 8'b11000100;
  assign _0521_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18302" *) 8'b11000101;
  assign _0522_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18364" *) 8'b11000110;
  assign _0523_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18426" *) 8'b11000111;
  assign _0524_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18488" *) 8'b11001000;
  assign _0525_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18550" *) 8'b11001001;
  assign _0526_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18612" *) 8'b11001010;
  assign _0527_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1866" *) reg2dp_lut_int_addr;
  assign _0528_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18674" *) 8'b11001011;
  assign _0529_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18736" *) 8'b11001100;
  assign _0530_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18798" *) 8'b11001101;
  assign _0531_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18860" *) 8'b11001110;
  assign _0532_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18922" *) 8'b11001111;
  assign _0533_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18984" *) 8'b11010000;
  assign _0534_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19046" *) 8'b11010001;
  assign _0535_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19108" *) 8'b11010010;
  assign _0536_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19170" *) 8'b11010011;
  assign _0537_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19232" *) 8'b11010100;
  assign _0538_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1928" *) 1'b1;
  assign _0539_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19294" *) 8'b11010101;
  assign _0540_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19356" *) 8'b11010110;
  assign _0541_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19418" *) 8'b11010111;
  assign _0542_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19480" *) 8'b11011000;
  assign _0543_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19542" *) 8'b11011001;
  assign _0544_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19604" *) 8'b11011010;
  assign _0545_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19666" *) 8'b11011011;
  assign _0546_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19728" *) 8'b11011100;
  assign _0547_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19790" *) 8'b11011101;
  assign _0548_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19852" *) 8'b11011110;
  assign _0549_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1990" *) 2'b10;
  assign _0550_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19914" *) 8'b11011111;
  assign _0551_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19976" *) 8'b11100000;
  assign _0552_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20038" *) 8'b11100001;
  assign _0553_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20100" *) 8'b11100010;
  assign _0554_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20162" *) 8'b11100011;
  assign _0555_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20224" *) 8'b11100100;
  assign _0556_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20286" *) 8'b11100101;
  assign _0557_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20348" *) 8'b11100110;
  assign _0558_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20410" *) 8'b11100111;
  assign _0559_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20472" *) 8'b11101000;
  assign _0560_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2052" *) 2'b11;
  assign _0561_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20534" *) 8'b11101001;
  assign _0562_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20596" *) 8'b11101010;
  assign _0563_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20658" *) 8'b11101011;
  assign _0564_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20720" *) 8'b11101100;
  assign _0565_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20782" *) 8'b11101101;
  assign _0566_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20844" *) 8'b11101110;
  assign _0567_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20906" *) 8'b11101111;
  assign _0568_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20968" *) 8'b11110000;
  assign _0569_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21030" *) 8'b11110001;
  assign _0570_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21092" *) 8'b11110010;
  assign _0571_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2114" *) 3'b100;
  assign _0572_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21154" *) 8'b11110011;
  assign _0573_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21216" *) 8'b11110100;
  assign _0574_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21278" *) 8'b11110101;
  assign _0575_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21340" *) 8'b11110110;
  assign _0576_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21402" *) 8'b11110111;
  assign _0577_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21464" *) 8'b11111000;
  assign _0578_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21526" *) 8'b11111001;
  assign _0579_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21588" *) 8'b11111010;
  assign _0580_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21650" *) 8'b11111011;
  assign _0581_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21712" *) 8'b11111100;
  assign _0582_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2176" *) 3'b101;
  assign _0583_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21774" *) 8'b11111101;
  assign _0584_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21836" *) 8'b11111110;
  assign _0585_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21898" *) 8'b11111111;
  assign _0586_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21960" *) 9'b100000000;
  assign _0587_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2238" *) 3'b110;
  assign _0588_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2300" *) 3'b111;
  assign _0589_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2362" *) 4'b1000;
  assign _0590_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2424" *) 4'b1001;
  assign _0591_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2486" *) 4'b1010;
  assign _0592_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2548" *) 4'b1011;
  assign _0593_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2610" *) 4'b1100;
  assign _0594_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2672" *) 4'b1101;
  assign _0595_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2734" *) 4'b1110;
  assign _0596_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2796" *) 4'b1111;
  assign _0597_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2858" *) 5'b10000;
  assign _0598_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2920" *) 5'b10001;
  assign _0599_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2982" *) 5'b10010;
  assign _0600_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3044" *) 5'b10011;
  assign _0601_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3106" *) 5'b10100;
  assign _0602_ = reg2dp_proc_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31126" *) 2'b10;
  assign _0603_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3168" *) 5'b10101;
  assign _0604_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3230" *) 5'b10110;
  assign _0605_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3292" *) 5'b10111;
  assign _0606_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3354" *) 5'b11000;
  assign _0607_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3416" *) 5'b11001;
  assign _0608_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3478" *) 5'b11010;
  assign _0609_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3540" *) 5'b11011;
  assign _0610_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3602" *) 5'b11100;
  assign _0611_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3664" *) 5'b11101;
  assign _0612_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3726" *) 5'b11110;
  assign _0613_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3788" *) 5'b11111;
  assign _0614_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3850" *) 6'b100000;
  assign _0615_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3912" *) 6'b100001;
  assign _0616_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3974" *) 6'b100010;
  assign _0617_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4036" *) 6'b100011;
  assign _0618_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4098" *) 6'b100100;
  assign _0619_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4160" *) 6'b100101;
  assign _0620_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4222" *) 6'b100110;
  assign _0621_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4284" *) 6'b100111;
  assign _0622_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4346" *) 6'b101000;
  assign _0623_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4408" *) 6'b101001;
  assign _0624_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4470" *) 6'b101010;
  assign _0625_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4532" *) 6'b101011;
  assign _0626_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4594" *) 6'b101100;
  assign _0627_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4656" *) 6'b101101;
  assign _0628_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4718" *) 6'b101110;
  assign _0629_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4780" *) 6'b101111;
  assign _0630_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4842" *) 6'b110000;
  assign _0631_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4904" *) 6'b110001;
  assign _0632_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4966" *) 6'b110010;
  assign _0633_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5028" *) 6'b110011;
  assign _0634_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5090" *) 6'b110100;
  assign _0635_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5152" *) 6'b110101;
  assign _0636_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5214" *) 6'b110110;
  assign _0637_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5276" *) 6'b110111;
  assign _0638_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5338" *) 6'b111000;
  assign _0639_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5400" *) 6'b111001;
  assign _0640_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5462" *) 6'b111010;
  assign _0641_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5524" *) 6'b111011;
  assign _0642_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5586" *) 6'b111100;
  assign _0643_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5648" *) 6'b111101;
  assign _0644_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5710" *) 6'b111110;
  assign _0645_ = reg2dp_lut_int_addr == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5772" *) 6'b111111;
  assign _0646_ = p1_pipe_ready_bc && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22230" *) idx2lut_pvld;
  assign _0647_ = dat_fifo_rd_prdy && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31594" *) dat_fifo_rd_pvld;
  assign _0648_ = p2_pipe_valid && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31609" *) p2_pipe_ready;
  assign p2_skid_catch = _0648_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31609" *) _0651_;
  assign _0649_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22219" *) p1_pipe_valid;
  assign lut_in_hybrid0 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22466" *) _0653_;
  assign lut_in_hybrid1 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22467" *) _0654_;
  assign lut_in_hybrid2 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22468" *) _0655_;
  assign lut_in_hybrid3 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22469" *) _0656_;
  assign _0650_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31583" *) p2_pipe_valid;
  assign _0651_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31609" *) lut2inp_prdy;
  assign _0652_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31610" *) p2_skid_catch;
  assign p1_pipe_ready_bc = cmd_fifo_wr_prdy || (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22219" *) _0649_;
  assign dat_fifo_rd_prdy = p2_pipe_ready || (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31583" *) _0650_;
  assign perf_lut_oflow_adv = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22389" *) perf_lut_oflow_add;
  assign perf_lut_uflow_adv = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22432" *) perf_lut_uflow_add;
  assign perf_lut_hybrid_adv = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22479" *) perf_lut_hybrid_add;
  assign perf_lut_le_hit_adv = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22522" *) perf_lut_le_hit_add;
  assign perf_lut_lo_hit_adv = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22565" *) perf_lut_lo_hit_add;
  assign _0653_ = p1_pipe_data[268] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22466" *) p1_pipe_data[272];
  assign _0654_ = p1_pipe_data[269] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22467" *) p1_pipe_data[273];
  assign _0655_ = p1_pipe_data[270] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22468" *) p1_pipe_data[274];
  assign _0656_ = p1_pipe_data[271] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22469" *) p1_pipe_data[275];
  assign out_flow0 = cmd_fifo_rd_pd[272] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31096" *) cmd_fifo_rd_pd[268];
  assign out_flow1 = cmd_fifo_rd_pd[273] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31097" *) cmd_fifo_rd_pd[269];
  assign out_flow2 = cmd_fifo_rd_pd[274] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31098" *) cmd_fifo_rd_pd[270];
  assign out_flow3 = cmd_fifo_rd_pd[275] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31099" *) cmd_fifo_rd_pd[271];
  always @(posedge nvdla_core_clk)
      p2_skid_data <= _0327_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      p2_pipe_ready <= 1'b1;
    else
      p2_pipe_ready <= p2_skid_ready;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      p2_skid_valid <= 1'b0;
    else
      p2_skid_valid <= _0328_;
  always @(posedge nvdla_core_clk)
      p2_pipe_data <= _0325_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      p2_pipe_valid <= 1'b0;
    else
      p2_pipe_valid <= _0326_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      perf_lut_lo_hit_cnt_cur <= 32'd0;
    else
      perf_lut_lo_hit_cnt_cur <= _0331_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      perf_lut_le_hit_cnt_cur <= 32'd0;
    else
      perf_lut_le_hit_cnt_cur <= _0330_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      perf_lut_hybrid_cnt_cur <= 32'd0;
    else
      perf_lut_hybrid_cnt_cur <= _0329_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      perf_lut_uflow_cnt_cur <= 32'd0;
    else
      perf_lut_uflow_cnt_cur <= _0333_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      perf_lut_oflow_cnt_cur <= 32'd0;
    else
      perf_lut_oflow_cnt_cur <= _0332_;
  always @(posedge nvdla_core_clk)
      p1_pipe_data <= _0323_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      p1_pipe_valid <= 1'b0;
    else
      p1_pipe_valid <= _0324_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_256 <= 16'b0000000000000000;
    else
      REG_lo_256 <= _0238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_255 <= 16'b0000000000000000;
    else
      REG_lo_255 <= _0237_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_254 <= 16'b0000000000000000;
    else
      REG_lo_254 <= _0236_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_253 <= 16'b0000000000000000;
    else
      REG_lo_253 <= _0235_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_252 <= 16'b0000000000000000;
    else
      REG_lo_252 <= _0234_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_251 <= 16'b0000000000000000;
    else
      REG_lo_251 <= _0233_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_250 <= 16'b0000000000000000;
    else
      REG_lo_250 <= _0232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_249 <= 16'b0000000000000000;
    else
      REG_lo_249 <= _0230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_248 <= 16'b0000000000000000;
    else
      REG_lo_248 <= _0229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_247 <= 16'b0000000000000000;
    else
      REG_lo_247 <= _0228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_246 <= 16'b0000000000000000;
    else
      REG_lo_246 <= _0227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_245 <= 16'b0000000000000000;
    else
      REG_lo_245 <= _0226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_244 <= 16'b0000000000000000;
    else
      REG_lo_244 <= _0225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_243 <= 16'b0000000000000000;
    else
      REG_lo_243 <= _0224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_242 <= 16'b0000000000000000;
    else
      REG_lo_242 <= _0223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_241 <= 16'b0000000000000000;
    else
      REG_lo_241 <= _0222_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_240 <= 16'b0000000000000000;
    else
      REG_lo_240 <= _0221_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_239 <= 16'b0000000000000000;
    else
      REG_lo_239 <= _0219_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_238 <= 16'b0000000000000000;
    else
      REG_lo_238 <= _0218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_237 <= 16'b0000000000000000;
    else
      REG_lo_237 <= _0217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_236 <= 16'b0000000000000000;
    else
      REG_lo_236 <= _0216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_235 <= 16'b0000000000000000;
    else
      REG_lo_235 <= _0215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_234 <= 16'b0000000000000000;
    else
      REG_lo_234 <= _0214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_233 <= 16'b0000000000000000;
    else
      REG_lo_233 <= _0213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_232 <= 16'b0000000000000000;
    else
      REG_lo_232 <= _0212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_231 <= 16'b0000000000000000;
    else
      REG_lo_231 <= _0211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_230 <= 16'b0000000000000000;
    else
      REG_lo_230 <= _0210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_229 <= 16'b0000000000000000;
    else
      REG_lo_229 <= _0208_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_228 <= 16'b0000000000000000;
    else
      REG_lo_228 <= _0207_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_227 <= 16'b0000000000000000;
    else
      REG_lo_227 <= _0206_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_226 <= 16'b0000000000000000;
    else
      REG_lo_226 <= _0205_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_225 <= 16'b0000000000000000;
    else
      REG_lo_225 <= _0204_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_224 <= 16'b0000000000000000;
    else
      REG_lo_224 <= _0203_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_223 <= 16'b0000000000000000;
    else
      REG_lo_223 <= _0202_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_222 <= 16'b0000000000000000;
    else
      REG_lo_222 <= _0201_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_221 <= 16'b0000000000000000;
    else
      REG_lo_221 <= _0200_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_220 <= 16'b0000000000000000;
    else
      REG_lo_220 <= _0199_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_219 <= 16'b0000000000000000;
    else
      REG_lo_219 <= _0197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_218 <= 16'b0000000000000000;
    else
      REG_lo_218 <= _0196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_217 <= 16'b0000000000000000;
    else
      REG_lo_217 <= _0195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_216 <= 16'b0000000000000000;
    else
      REG_lo_216 <= _0194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_215 <= 16'b0000000000000000;
    else
      REG_lo_215 <= _0193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_214 <= 16'b0000000000000000;
    else
      REG_lo_214 <= _0192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_213 <= 16'b0000000000000000;
    else
      REG_lo_213 <= _0191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_212 <= 16'b0000000000000000;
    else
      REG_lo_212 <= _0190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_211 <= 16'b0000000000000000;
    else
      REG_lo_211 <= _0189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_210 <= 16'b0000000000000000;
    else
      REG_lo_210 <= _0188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_209 <= 16'b0000000000000000;
    else
      REG_lo_209 <= _0186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_208 <= 16'b0000000000000000;
    else
      REG_lo_208 <= _0185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_207 <= 16'b0000000000000000;
    else
      REG_lo_207 <= _0184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_206 <= 16'b0000000000000000;
    else
      REG_lo_206 <= _0183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_205 <= 16'b0000000000000000;
    else
      REG_lo_205 <= _0182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_204 <= 16'b0000000000000000;
    else
      REG_lo_204 <= _0181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_203 <= 16'b0000000000000000;
    else
      REG_lo_203 <= _0180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_202 <= 16'b0000000000000000;
    else
      REG_lo_202 <= _0179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_201 <= 16'b0000000000000000;
    else
      REG_lo_201 <= _0178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_200 <= 16'b0000000000000000;
    else
      REG_lo_200 <= _0177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_199 <= 16'b0000000000000000;
    else
      REG_lo_199 <= _0174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_198 <= 16'b0000000000000000;
    else
      REG_lo_198 <= _0173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_197 <= 16'b0000000000000000;
    else
      REG_lo_197 <= _0172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_196 <= 16'b0000000000000000;
    else
      REG_lo_196 <= _0171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_195 <= 16'b0000000000000000;
    else
      REG_lo_195 <= _0170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_194 <= 16'b0000000000000000;
    else
      REG_lo_194 <= _0169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_193 <= 16'b0000000000000000;
    else
      REG_lo_193 <= _0168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_192 <= 16'b0000000000000000;
    else
      REG_lo_192 <= _0167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_191 <= 16'b0000000000000000;
    else
      REG_lo_191 <= _0166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_190 <= 16'b0000000000000000;
    else
      REG_lo_190 <= _0165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_189 <= 16'b0000000000000000;
    else
      REG_lo_189 <= _0163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_188 <= 16'b0000000000000000;
    else
      REG_lo_188 <= _0162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_187 <= 16'b0000000000000000;
    else
      REG_lo_187 <= _0161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_186 <= 16'b0000000000000000;
    else
      REG_lo_186 <= _0160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_185 <= 16'b0000000000000000;
    else
      REG_lo_185 <= _0159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_184 <= 16'b0000000000000000;
    else
      REG_lo_184 <= _0158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_183 <= 16'b0000000000000000;
    else
      REG_lo_183 <= _0157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_182 <= 16'b0000000000000000;
    else
      REG_lo_182 <= _0156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_181 <= 16'b0000000000000000;
    else
      REG_lo_181 <= _0155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_180 <= 16'b0000000000000000;
    else
      REG_lo_180 <= _0154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_179 <= 16'b0000000000000000;
    else
      REG_lo_179 <= _0152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_178 <= 16'b0000000000000000;
    else
      REG_lo_178 <= _0151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_177 <= 16'b0000000000000000;
    else
      REG_lo_177 <= _0150_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_176 <= 16'b0000000000000000;
    else
      REG_lo_176 <= _0149_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_175 <= 16'b0000000000000000;
    else
      REG_lo_175 <= _0148_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_174 <= 16'b0000000000000000;
    else
      REG_lo_174 <= _0147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_173 <= 16'b0000000000000000;
    else
      REG_lo_173 <= _0146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_172 <= 16'b0000000000000000;
    else
      REG_lo_172 <= _0145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_171 <= 16'b0000000000000000;
    else
      REG_lo_171 <= _0144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_170 <= 16'b0000000000000000;
    else
      REG_lo_170 <= _0143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_169 <= 16'b0000000000000000;
    else
      REG_lo_169 <= _0141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_168 <= 16'b0000000000000000;
    else
      REG_lo_168 <= _0140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_167 <= 16'b0000000000000000;
    else
      REG_lo_167 <= _0139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_166 <= 16'b0000000000000000;
    else
      REG_lo_166 <= _0138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_165 <= 16'b0000000000000000;
    else
      REG_lo_165 <= _0137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_164 <= 16'b0000000000000000;
    else
      REG_lo_164 <= _0136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_163 <= 16'b0000000000000000;
    else
      REG_lo_163 <= _0135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_162 <= 16'b0000000000000000;
    else
      REG_lo_162 <= _0134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_161 <= 16'b0000000000000000;
    else
      REG_lo_161 <= _0133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_160 <= 16'b0000000000000000;
    else
      REG_lo_160 <= _0132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_159 <= 16'b0000000000000000;
    else
      REG_lo_159 <= _0130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_158 <= 16'b0000000000000000;
    else
      REG_lo_158 <= _0129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_157 <= 16'b0000000000000000;
    else
      REG_lo_157 <= _0128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_156 <= 16'b0000000000000000;
    else
      REG_lo_156 <= _0127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_155 <= 16'b0000000000000000;
    else
      REG_lo_155 <= _0126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_154 <= 16'b0000000000000000;
    else
      REG_lo_154 <= _0125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_153 <= 16'b0000000000000000;
    else
      REG_lo_153 <= _0124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_152 <= 16'b0000000000000000;
    else
      REG_lo_152 <= _0123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_151 <= 16'b0000000000000000;
    else
      REG_lo_151 <= _0122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_150 <= 16'b0000000000000000;
    else
      REG_lo_150 <= _0121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_149 <= 16'b0000000000000000;
    else
      REG_lo_149 <= _0119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_148 <= 16'b0000000000000000;
    else
      REG_lo_148 <= _0118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_147 <= 16'b0000000000000000;
    else
      REG_lo_147 <= _0117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_146 <= 16'b0000000000000000;
    else
      REG_lo_146 <= _0116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_145 <= 16'b0000000000000000;
    else
      REG_lo_145 <= _0115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_144 <= 16'b0000000000000000;
    else
      REG_lo_144 <= _0114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_143 <= 16'b0000000000000000;
    else
      REG_lo_143 <= _0113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_142 <= 16'b0000000000000000;
    else
      REG_lo_142 <= _0112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_141 <= 16'b0000000000000000;
    else
      REG_lo_141 <= _0111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_140 <= 16'b0000000000000000;
    else
      REG_lo_140 <= _0110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_139 <= 16'b0000000000000000;
    else
      REG_lo_139 <= _0108_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_138 <= 16'b0000000000000000;
    else
      REG_lo_138 <= _0107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_137 <= 16'b0000000000000000;
    else
      REG_lo_137 <= _0106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_136 <= 16'b0000000000000000;
    else
      REG_lo_136 <= _0105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_135 <= 16'b0000000000000000;
    else
      REG_lo_135 <= _0104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_134 <= 16'b0000000000000000;
    else
      REG_lo_134 <= _0103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_133 <= 16'b0000000000000000;
    else
      REG_lo_133 <= _0102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_132 <= 16'b0000000000000000;
    else
      REG_lo_132 <= _0101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_131 <= 16'b0000000000000000;
    else
      REG_lo_131 <= _0100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_130 <= 16'b0000000000000000;
    else
      REG_lo_130 <= _0099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_129 <= 16'b0000000000000000;
    else
      REG_lo_129 <= _0097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_128 <= 16'b0000000000000000;
    else
      REG_lo_128 <= _0096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_127 <= 16'b0000000000000000;
    else
      REG_lo_127 <= _0095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_126 <= 16'b0000000000000000;
    else
      REG_lo_126 <= _0094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_125 <= 16'b0000000000000000;
    else
      REG_lo_125 <= _0093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_124 <= 16'b0000000000000000;
    else
      REG_lo_124 <= _0092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_123 <= 16'b0000000000000000;
    else
      REG_lo_123 <= _0091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_122 <= 16'b0000000000000000;
    else
      REG_lo_122 <= _0090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_121 <= 16'b0000000000000000;
    else
      REG_lo_121 <= _0089_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_120 <= 16'b0000000000000000;
    else
      REG_lo_120 <= _0088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_119 <= 16'b0000000000000000;
    else
      REG_lo_119 <= _0086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_118 <= 16'b0000000000000000;
    else
      REG_lo_118 <= _0085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_117 <= 16'b0000000000000000;
    else
      REG_lo_117 <= _0084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_116 <= 16'b0000000000000000;
    else
      REG_lo_116 <= _0083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_115 <= 16'b0000000000000000;
    else
      REG_lo_115 <= _0082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_114 <= 16'b0000000000000000;
    else
      REG_lo_114 <= _0081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_113 <= 16'b0000000000000000;
    else
      REG_lo_113 <= _0080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_112 <= 16'b0000000000000000;
    else
      REG_lo_112 <= _0079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_111 <= 16'b0000000000000000;
    else
      REG_lo_111 <= _0078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_110 <= 16'b0000000000000000;
    else
      REG_lo_110 <= _0077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_109 <= 16'b0000000000000000;
    else
      REG_lo_109 <= _0075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_108 <= 16'b0000000000000000;
    else
      REG_lo_108 <= _0074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_107 <= 16'b0000000000000000;
    else
      REG_lo_107 <= _0073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_106 <= 16'b0000000000000000;
    else
      REG_lo_106 <= _0072_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_105 <= 16'b0000000000000000;
    else
      REG_lo_105 <= _0071_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_104 <= 16'b0000000000000000;
    else
      REG_lo_104 <= _0070_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_103 <= 16'b0000000000000000;
    else
      REG_lo_103 <= _0069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_102 <= 16'b0000000000000000;
    else
      REG_lo_102 <= _0068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_101 <= 16'b0000000000000000;
    else
      REG_lo_101 <= _0067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_100 <= 16'b0000000000000000;
    else
      REG_lo_100 <= _0066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_99 <= 16'b0000000000000000;
    else
      REG_lo_99 <= _0320_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_98 <= 16'b0000000000000000;
    else
      REG_lo_98 <= _0319_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_97 <= 16'b0000000000000000;
    else
      REG_lo_97 <= _0318_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_96 <= 16'b0000000000000000;
    else
      REG_lo_96 <= _0317_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_95 <= 16'b0000000000000000;
    else
      REG_lo_95 <= _0316_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_94 <= 16'b0000000000000000;
    else
      REG_lo_94 <= _0315_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_93 <= 16'b0000000000000000;
    else
      REG_lo_93 <= _0314_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_92 <= 16'b0000000000000000;
    else
      REG_lo_92 <= _0313_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_91 <= 16'b0000000000000000;
    else
      REG_lo_91 <= _0312_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_90 <= 16'b0000000000000000;
    else
      REG_lo_90 <= _0311_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_89 <= 16'b0000000000000000;
    else
      REG_lo_89 <= _0309_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_88 <= 16'b0000000000000000;
    else
      REG_lo_88 <= _0308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_87 <= 16'b0000000000000000;
    else
      REG_lo_87 <= _0307_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_86 <= 16'b0000000000000000;
    else
      REG_lo_86 <= _0306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_85 <= 16'b0000000000000000;
    else
      REG_lo_85 <= _0305_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_84 <= 16'b0000000000000000;
    else
      REG_lo_84 <= _0304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_83 <= 16'b0000000000000000;
    else
      REG_lo_83 <= _0303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_82 <= 16'b0000000000000000;
    else
      REG_lo_82 <= _0302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_81 <= 16'b0000000000000000;
    else
      REG_lo_81 <= _0301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_80 <= 16'b0000000000000000;
    else
      REG_lo_80 <= _0300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_79 <= 16'b0000000000000000;
    else
      REG_lo_79 <= _0298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_78 <= 16'b0000000000000000;
    else
      REG_lo_78 <= _0297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_77 <= 16'b0000000000000000;
    else
      REG_lo_77 <= _0296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_76 <= 16'b0000000000000000;
    else
      REG_lo_76 <= _0295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_75 <= 16'b0000000000000000;
    else
      REG_lo_75 <= _0294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_74 <= 16'b0000000000000000;
    else
      REG_lo_74 <= _0293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_73 <= 16'b0000000000000000;
    else
      REG_lo_73 <= _0292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_72 <= 16'b0000000000000000;
    else
      REG_lo_72 <= _0291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_71 <= 16'b0000000000000000;
    else
      REG_lo_71 <= _0290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_70 <= 16'b0000000000000000;
    else
      REG_lo_70 <= _0289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_69 <= 16'b0000000000000000;
    else
      REG_lo_69 <= _0287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_68 <= 16'b0000000000000000;
    else
      REG_lo_68 <= _0286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_67 <= 16'b0000000000000000;
    else
      REG_lo_67 <= _0285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_66 <= 16'b0000000000000000;
    else
      REG_lo_66 <= _0284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_65 <= 16'b0000000000000000;
    else
      REG_lo_65 <= _0283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_64 <= 16'b0000000000000000;
    else
      REG_lo_64 <= _0282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_63 <= 16'b0000000000000000;
    else
      REG_lo_63 <= _0281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_62 <= 16'b0000000000000000;
    else
      REG_lo_62 <= _0280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_61 <= 16'b0000000000000000;
    else
      REG_lo_61 <= _0279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_60 <= 16'b0000000000000000;
    else
      REG_lo_60 <= _0278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_59 <= 16'b0000000000000000;
    else
      REG_lo_59 <= _0276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_58 <= 16'b0000000000000000;
    else
      REG_lo_58 <= _0275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_57 <= 16'b0000000000000000;
    else
      REG_lo_57 <= _0274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_56 <= 16'b0000000000000000;
    else
      REG_lo_56 <= _0273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_55 <= 16'b0000000000000000;
    else
      REG_lo_55 <= _0272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_54 <= 16'b0000000000000000;
    else
      REG_lo_54 <= _0271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_53 <= 16'b0000000000000000;
    else
      REG_lo_53 <= _0270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_52 <= 16'b0000000000000000;
    else
      REG_lo_52 <= _0269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_51 <= 16'b0000000000000000;
    else
      REG_lo_51 <= _0268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_50 <= 16'b0000000000000000;
    else
      REG_lo_50 <= _0267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_49 <= 16'b0000000000000000;
    else
      REG_lo_49 <= _0265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_48 <= 16'b0000000000000000;
    else
      REG_lo_48 <= _0264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_47 <= 16'b0000000000000000;
    else
      REG_lo_47 <= _0263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_46 <= 16'b0000000000000000;
    else
      REG_lo_46 <= _0262_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_45 <= 16'b0000000000000000;
    else
      REG_lo_45 <= _0261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_44 <= 16'b0000000000000000;
    else
      REG_lo_44 <= _0260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_43 <= 16'b0000000000000000;
    else
      REG_lo_43 <= _0259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_42 <= 16'b0000000000000000;
    else
      REG_lo_42 <= _0258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_41 <= 16'b0000000000000000;
    else
      REG_lo_41 <= _0257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_40 <= 16'b0000000000000000;
    else
      REG_lo_40 <= _0256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_39 <= 16'b0000000000000000;
    else
      REG_lo_39 <= _0254_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_38 <= 16'b0000000000000000;
    else
      REG_lo_38 <= _0253_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_37 <= 16'b0000000000000000;
    else
      REG_lo_37 <= _0252_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_36 <= 16'b0000000000000000;
    else
      REG_lo_36 <= _0251_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_35 <= 16'b0000000000000000;
    else
      REG_lo_35 <= _0250_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_34 <= 16'b0000000000000000;
    else
      REG_lo_34 <= _0249_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_33 <= 16'b0000000000000000;
    else
      REG_lo_33 <= _0248_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_32 <= 16'b0000000000000000;
    else
      REG_lo_32 <= _0247_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_31 <= 16'b0000000000000000;
    else
      REG_lo_31 <= _0246_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_30 <= 16'b0000000000000000;
    else
      REG_lo_30 <= _0245_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_29 <= 16'b0000000000000000;
    else
      REG_lo_29 <= _0243_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_28 <= 16'b0000000000000000;
    else
      REG_lo_28 <= _0242_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_27 <= 16'b0000000000000000;
    else
      REG_lo_27 <= _0241_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_26 <= 16'b0000000000000000;
    else
      REG_lo_26 <= _0240_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_25 <= 16'b0000000000000000;
    else
      REG_lo_25 <= _0239_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_24 <= 16'b0000000000000000;
    else
      REG_lo_24 <= _0231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_23 <= 16'b0000000000000000;
    else
      REG_lo_23 <= _0220_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_22 <= 16'b0000000000000000;
    else
      REG_lo_22 <= _0209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_21 <= 16'b0000000000000000;
    else
      REG_lo_21 <= _0198_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_20 <= 16'b0000000000000000;
    else
      REG_lo_20 <= _0187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_19 <= 16'b0000000000000000;
    else
      REG_lo_19 <= _0175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_18 <= 16'b0000000000000000;
    else
      REG_lo_18 <= _0164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_17 <= 16'b0000000000000000;
    else
      REG_lo_17 <= _0153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_16 <= 16'b0000000000000000;
    else
      REG_lo_16 <= _0142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_15 <= 16'b0000000000000000;
    else
      REG_lo_15 <= _0131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_14 <= 16'b0000000000000000;
    else
      REG_lo_14 <= _0120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_13 <= 16'b0000000000000000;
    else
      REG_lo_13 <= _0109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_12 <= 16'b0000000000000000;
    else
      REG_lo_12 <= _0098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_11 <= 16'b0000000000000000;
    else
      REG_lo_11 <= _0087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_10 <= 16'b0000000000000000;
    else
      REG_lo_10 <= _0076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_9 <= 16'b0000000000000000;
    else
      REG_lo_9 <= _0321_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_8 <= 16'b0000000000000000;
    else
      REG_lo_8 <= _0310_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_7 <= 16'b0000000000000000;
    else
      REG_lo_7 <= _0299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_6 <= 16'b0000000000000000;
    else
      REG_lo_6 <= _0288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_5 <= 16'b0000000000000000;
    else
      REG_lo_5 <= _0277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_4 <= 16'b0000000000000000;
    else
      REG_lo_4 <= _0266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_3 <= 16'b0000000000000000;
    else
      REG_lo_3 <= _0255_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_2 <= 16'b0000000000000000;
    else
      REG_lo_2 <= _0244_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_1 <= 16'b0000000000000000;
    else
      REG_lo_1 <= _0176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_lo_0 <= 16'b0000000000000000;
    else
      REG_lo_0 <= _0065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_64 <= 16'b0000000000000000;
    else
      REG_le_64 <= _0060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_63 <= 16'b0000000000000000;
    else
      REG_le_63 <= _0059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_62 <= 16'b0000000000000000;
    else
      REG_le_62 <= _0058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_61 <= 16'b0000000000000000;
    else
      REG_le_61 <= _0057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_60 <= 16'b0000000000000000;
    else
      REG_le_60 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_59 <= 16'b0000000000000000;
    else
      REG_le_59 <= _0054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_58 <= 16'b0000000000000000;
    else
      REG_le_58 <= _0053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_57 <= 16'b0000000000000000;
    else
      REG_le_57 <= _0052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_56 <= 16'b0000000000000000;
    else
      REG_le_56 <= _0051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_55 <= 16'b0000000000000000;
    else
      REG_le_55 <= _0050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_54 <= 16'b0000000000000000;
    else
      REG_le_54 <= _0049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_53 <= 16'b0000000000000000;
    else
      REG_le_53 <= _0048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_52 <= 16'b0000000000000000;
    else
      REG_le_52 <= _0047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_51 <= 16'b0000000000000000;
    else
      REG_le_51 <= _0046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_50 <= 16'b0000000000000000;
    else
      REG_le_50 <= _0045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_49 <= 16'b0000000000000000;
    else
      REG_le_49 <= _0043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_48 <= 16'b0000000000000000;
    else
      REG_le_48 <= _0042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_47 <= 16'b0000000000000000;
    else
      REG_le_47 <= _0041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_46 <= 16'b0000000000000000;
    else
      REG_le_46 <= _0040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_45 <= 16'b0000000000000000;
    else
      REG_le_45 <= _0039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_44 <= 16'b0000000000000000;
    else
      REG_le_44 <= _0038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_43 <= 16'b0000000000000000;
    else
      REG_le_43 <= _0037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_42 <= 16'b0000000000000000;
    else
      REG_le_42 <= _0036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_41 <= 16'b0000000000000000;
    else
      REG_le_41 <= _0035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_40 <= 16'b0000000000000000;
    else
      REG_le_40 <= _0034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_39 <= 16'b0000000000000000;
    else
      REG_le_39 <= _0032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_38 <= 16'b0000000000000000;
    else
      REG_le_38 <= _0031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_37 <= 16'b0000000000000000;
    else
      REG_le_37 <= _0030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_36 <= 16'b0000000000000000;
    else
      REG_le_36 <= _0029_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_35 <= 16'b0000000000000000;
    else
      REG_le_35 <= _0028_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_34 <= 16'b0000000000000000;
    else
      REG_le_34 <= _0027_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_33 <= 16'b0000000000000000;
    else
      REG_le_33 <= _0026_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_32 <= 16'b0000000000000000;
    else
      REG_le_32 <= _0025_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_31 <= 16'b0000000000000000;
    else
      REG_le_31 <= _0024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_30 <= 16'b0000000000000000;
    else
      REG_le_30 <= _0023_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_29 <= 16'b0000000000000000;
    else
      REG_le_29 <= _0021_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_28 <= 16'b0000000000000000;
    else
      REG_le_28 <= _0020_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_27 <= 16'b0000000000000000;
    else
      REG_le_27 <= _0019_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_26 <= 16'b0000000000000000;
    else
      REG_le_26 <= _0018_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_25 <= 16'b0000000000000000;
    else
      REG_le_25 <= _0017_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_24 <= 16'b0000000000000000;
    else
      REG_le_24 <= _0016_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_23 <= 16'b0000000000000000;
    else
      REG_le_23 <= _0015_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_22 <= 16'b0000000000000000;
    else
      REG_le_22 <= _0014_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_21 <= 16'b0000000000000000;
    else
      REG_le_21 <= _0013_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_20 <= 16'b0000000000000000;
    else
      REG_le_20 <= _0012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_19 <= 16'b0000000000000000;
    else
      REG_le_19 <= _0010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_18 <= 16'b0000000000000000;
    else
      REG_le_18 <= _0009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_17 <= 16'b0000000000000000;
    else
      REG_le_17 <= _0008_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_16 <= 16'b0000000000000000;
    else
      REG_le_16 <= _0007_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_15 <= 16'b0000000000000000;
    else
      REG_le_15 <= _0006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_14 <= 16'b0000000000000000;
    else
      REG_le_14 <= _0005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_13 <= 16'b0000000000000000;
    else
      REG_le_13 <= _0004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_12 <= 16'b0000000000000000;
    else
      REG_le_12 <= _0003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_11 <= 16'b0000000000000000;
    else
      REG_le_11 <= _0002_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_10 <= 16'b0000000000000000;
    else
      REG_le_10 <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_9 <= 16'b0000000000000000;
    else
      REG_le_9 <= _0064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_8 <= 16'b0000000000000000;
    else
      REG_le_8 <= _0063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_7 <= 16'b0000000000000000;
    else
      REG_le_7 <= _0062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_6 <= 16'b0000000000000000;
    else
      REG_le_6 <= _0061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_5 <= 16'b0000000000000000;
    else
      REG_le_5 <= _0055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_4 <= 16'b0000000000000000;
    else
      REG_le_4 <= _0044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_3 <= 16'b0000000000000000;
    else
      REG_le_3 <= _0033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_2 <= 16'b0000000000000000;
    else
      REG_le_2 <= _0022_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_1 <= 16'b0000000000000000;
    else
      REG_le_1 <= _0011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      REG_le_0 <= 16'b0000000000000000;
    else
      REG_le_0 <= _0000_;
  assign _0367_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31330" *) reg2dp_lut_lo_end : reg2dp_lut_le_end;
  assign _0375_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31330" *) reg2dp_lut_lo_slope_oflow_shift : reg2dp_lut_le_slope_oflow_shift;
  assign _0371_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31330" *) reg2dp_lut_lo_slope_oflow_scale : reg2dp_lut_le_slope_oflow_scale;
  assign _0362_ = cmd_fifo_rd_pd[271] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31329" *) _0375_ : 5'b00000;
  assign _0358_ = cmd_fifo_rd_pd[271] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31329" *) _0371_ : 16'b0000000000000000;
  assign _0354_ = cmd_fifo_rd_pd[271] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31329" *) _0367_ : 32'd0;
  assign _0363_ = _0602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31312" *) { 1'b0, _0322_, 23'b00000000000000000000000 } : _2715_;
  assign _0350_ = reg2dp_lut_le_function ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31311" *) 32'd0 : _0363_;
  assign _0337_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31307" *) 32'd0 : _0350_;
  assign _0341_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31307" *) reg2dp_lut_lo_start : reg2dp_lut_le_start;
  assign _0349_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31307" *) reg2dp_lut_lo_slope_uflow_shift : reg2dp_lut_le_slope_uflow_shift;
  assign _0345_ = cmd_fifo_rd_pd[279] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31307" *) reg2dp_lut_lo_slope_uflow_scale : reg2dp_lut_le_slope_uflow_scale;
  assign out_shift3 = cmd_fifo_rd_pd[275] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31306" *) _0349_ : _0362_;
  assign out_scale3 = cmd_fifo_rd_pd[275] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31306" *) _0345_ : _0358_;
  assign out_offset3 = cmd_fifo_rd_pd[275] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31306" *) _0341_ : _0354_;
  assign out_bias3 = cmd_fifo_rd_pd[275] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31306" *) _0337_ : 32'd0;
  assign _0366_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31268" *) reg2dp_lut_lo_end : reg2dp_lut_le_end;
  assign _0374_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31268" *) reg2dp_lut_lo_slope_oflow_shift : reg2dp_lut_le_slope_oflow_shift;
  assign _0370_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31268" *) reg2dp_lut_lo_slope_oflow_scale : reg2dp_lut_le_slope_oflow_scale;
  assign _0361_ = cmd_fifo_rd_pd[270] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31267" *) _0374_ : 5'b00000;
  assign _0357_ = cmd_fifo_rd_pd[270] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31267" *) _0370_ : 16'b0000000000000000;
  assign _0353_ = cmd_fifo_rd_pd[270] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31267" *) _0366_ : 32'd0;
  assign _0336_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31245" *) 32'd0 : _0350_;
  assign _0340_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31245" *) reg2dp_lut_lo_start : reg2dp_lut_le_start;
  assign _0348_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31245" *) reg2dp_lut_lo_slope_uflow_shift : reg2dp_lut_le_slope_uflow_shift;
  assign _0344_ = cmd_fifo_rd_pd[278] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31245" *) reg2dp_lut_lo_slope_uflow_scale : reg2dp_lut_le_slope_uflow_scale;
  assign out_shift2 = cmd_fifo_rd_pd[274] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31244" *) _0348_ : _0361_;
  assign out_scale2 = cmd_fifo_rd_pd[274] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31244" *) _0344_ : _0357_;
  assign out_offset2 = cmd_fifo_rd_pd[274] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31244" *) _0340_ : _0353_;
  assign out_bias2 = cmd_fifo_rd_pd[274] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31244" *) _0336_ : 32'd0;
  assign _0365_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31206" *) reg2dp_lut_lo_end : reg2dp_lut_le_end;
  assign _0373_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31206" *) reg2dp_lut_lo_slope_oflow_shift : reg2dp_lut_le_slope_oflow_shift;
  assign _0369_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31206" *) reg2dp_lut_lo_slope_oflow_scale : reg2dp_lut_le_slope_oflow_scale;
  assign _0360_ = cmd_fifo_rd_pd[269] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31205" *) _0373_ : 5'b00000;
  assign _0356_ = cmd_fifo_rd_pd[269] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31205" *) _0369_ : 16'b0000000000000000;
  assign _0352_ = cmd_fifo_rd_pd[269] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31205" *) _0365_ : 32'd0;
  assign _0335_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31183" *) 32'd0 : _0350_;
  assign _0339_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31183" *) reg2dp_lut_lo_start : reg2dp_lut_le_start;
  assign _0347_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31183" *) reg2dp_lut_lo_slope_uflow_shift : reg2dp_lut_le_slope_uflow_shift;
  assign _0343_ = cmd_fifo_rd_pd[277] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31183" *) reg2dp_lut_lo_slope_uflow_scale : reg2dp_lut_le_slope_uflow_scale;
  assign out_shift1 = cmd_fifo_rd_pd[273] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31182" *) _0347_ : _0360_;
  assign out_scale1 = cmd_fifo_rd_pd[273] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31182" *) _0343_ : _0356_;
  assign out_offset1 = cmd_fifo_rd_pd[273] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31182" *) _0339_ : _0352_;
  assign out_bias1 = cmd_fifo_rd_pd[273] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31182" *) _0335_ : 32'd0;
  assign _0364_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31144" *) reg2dp_lut_lo_end : reg2dp_lut_le_end;
  assign _0372_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31144" *) reg2dp_lut_lo_slope_oflow_shift : reg2dp_lut_le_slope_oflow_shift;
  assign _0368_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31144" *) reg2dp_lut_lo_slope_oflow_scale : reg2dp_lut_le_slope_oflow_scale;
  assign _0359_ = cmd_fifo_rd_pd[268] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31143" *) _0372_ : 5'b00000;
  assign _0355_ = cmd_fifo_rd_pd[268] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31143" *) _0368_ : 16'b0000000000000000;
  assign _0351_ = cmd_fifo_rd_pd[268] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31143" *) _0364_ : 32'd0;
  assign _0334_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31121" *) 32'd0 : _0350_;
  assign _0338_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31121" *) reg2dp_lut_lo_start : reg2dp_lut_le_start;
  assign _0346_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31121" *) reg2dp_lut_lo_slope_uflow_shift : reg2dp_lut_le_slope_uflow_shift;
  assign _0342_ = cmd_fifo_rd_pd[276] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31121" *) reg2dp_lut_lo_slope_uflow_scale : reg2dp_lut_le_slope_uflow_scale;
  assign out_shift0 = cmd_fifo_rd_pd[272] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31120" *) _0346_ : _0359_;
  assign out_scale0 = cmd_fifo_rd_pd[272] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31120" *) _0342_ : _0355_;
  assign out_offset0 = cmd_fifo_rd_pd[272] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31120" *) _0338_ : _0351_;
  assign out_bias0 = cmd_fifo_rd_pd[272] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31120" *) _0334_ : 32'd0;
  function [15:0] _3746_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30984|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _3746_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _3746_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _3746_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _3746_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _3746_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _3746_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _3746_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _3746_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _3746_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _3746_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _3746_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _3746_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _3746_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _3746_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _3746_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _3746_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _3746_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _3746_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _3746_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _3746_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _3746_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _3746_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _3746_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _3746_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _3746_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _3746_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _3746_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _3746_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _3746_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _3746_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _3746_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _3746_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _3746_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _3746_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _3746_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _3746_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _3746_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _3746_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _3746_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _3746_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _3746_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _3746_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _3746_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _3746_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _3746_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _3746_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _3746_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _3746_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _3746_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _3746_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _3746_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _3746_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _3746_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _3746_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _3746_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _3746_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _3746_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _3746_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _3746_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _3746_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _3746_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _3746_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _3746_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _3746_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _3746_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _3746_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _3746_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _3746_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _3746_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _3746_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _3746_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _3746_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _3746_ = b[4095:4080];
      default:
        _3746_ = a;
    endcase
  endfunction
  assign lo_data1_3 = _3746_(16'b0000000000000000, { REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_, _0774_, _0773_, _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0676_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0665_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_ });
  assign _0657_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30984|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 9'b100000000;
  assign _0658_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30983|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111111;
  assign _0659_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30982|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111110;
  assign _0660_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30981|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111101;
  assign _0661_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30980|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111100;
  assign _0662_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30979|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111011;
  assign _0663_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30978|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111010;
  assign _0664_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30977|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111001;
  assign _0665_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30976|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11111000;
  assign _0666_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30975|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110111;
  assign _0667_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30974|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110110;
  assign _0668_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30973|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110101;
  assign _0669_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30972|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110100;
  assign _0670_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30971|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110011;
  assign _0671_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30970|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110010;
  assign _0672_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30969|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110001;
  assign _0673_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30968|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11110000;
  assign _0674_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30967|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101111;
  assign _0675_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30966|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101110;
  assign _0676_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30965|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101101;
  assign _0677_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30964|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101100;
  assign _0678_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30963|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101011;
  assign _0679_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30962|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101010;
  assign _0680_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30961|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101001;
  assign _0681_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30960|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11101000;
  assign _0682_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30959|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100111;
  assign _0683_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30958|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100110;
  assign _0684_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30957|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100101;
  assign _0685_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30956|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100100;
  assign _0686_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30955|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100011;
  assign _0687_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30954|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100010;
  assign _0688_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30953|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100001;
  assign _0689_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30952|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11100000;
  assign _0690_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30951|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011111;
  assign _0691_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30950|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011110;
  assign _0692_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30949|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011101;
  assign _0693_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30948|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011100;
  assign _0694_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30947|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011011;
  assign _0695_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30946|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011010;
  assign _0696_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30945|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011001;
  assign _0697_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30944|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11011000;
  assign _0698_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30943|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010111;
  assign _0699_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30942|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010110;
  assign _0700_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30941|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010101;
  assign _0701_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30940|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010100;
  assign _0702_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30939|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010011;
  assign _0703_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30938|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010010;
  assign _0704_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30937|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010001;
  assign _0705_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30936|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11010000;
  assign _0706_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30935|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001111;
  assign _0707_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30934|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001110;
  assign _0708_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30933|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001101;
  assign _0709_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30932|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001100;
  assign _0710_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30931|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001011;
  assign _0711_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30930|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001010;
  assign _0712_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30929|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001001;
  assign _0713_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30928|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11001000;
  assign _0714_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30927|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000111;
  assign _0715_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30926|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000110;
  assign _0716_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30925|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000101;
  assign _0717_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30924|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000100;
  assign _0718_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30923|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000011;
  assign _0719_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30922|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000010;
  assign _0720_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30921|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000001;
  assign _0721_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30920|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b11000000;
  assign _0722_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30919|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111111;
  assign _0723_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30918|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111110;
  assign _0724_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30917|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111101;
  assign _0725_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30916|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111100;
  assign _0726_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30915|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111011;
  assign _0727_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30914|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111010;
  assign _0728_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30913|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111001;
  assign _0729_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30912|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10111000;
  assign _0730_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30911|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110111;
  assign _0731_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30910|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110110;
  assign _0732_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30909|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110101;
  assign _0733_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30908|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110100;
  assign _0734_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30907|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110011;
  assign _0735_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30906|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110010;
  assign _0736_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30905|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110001;
  assign _0737_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30904|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10110000;
  assign _0738_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30903|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101111;
  assign _0739_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30902|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101110;
  assign _0740_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30901|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101101;
  assign _0741_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30900|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101100;
  assign _0742_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30899|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101011;
  assign _0743_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30898|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101010;
  assign _0744_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30897|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101001;
  assign _0745_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30896|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10101000;
  assign _0746_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30895|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100111;
  assign _0747_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30894|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100110;
  assign _0748_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30893|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100101;
  assign _0749_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30892|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100100;
  assign _0750_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30891|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100011;
  assign _0751_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30890|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100010;
  assign _0752_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30889|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100001;
  assign _0753_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30888|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10100000;
  assign _0754_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30887|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011111;
  assign _0755_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30886|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011110;
  assign _0756_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30885|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011101;
  assign _0757_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30884|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011100;
  assign _0758_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30883|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011011;
  assign _0759_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30882|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011010;
  assign _0760_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30881|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011001;
  assign _0761_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30880|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10011000;
  assign _0762_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30879|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010111;
  assign _0763_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30878|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010110;
  assign _0764_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30877|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010101;
  assign _0765_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30876|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010100;
  assign _0766_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30875|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010011;
  assign _0767_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30874|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010010;
  assign _0768_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30873|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010001;
  assign _0769_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30872|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10010000;
  assign _0770_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30871|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001111;
  assign _0771_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30870|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001110;
  assign _0772_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30869|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001101;
  assign _0773_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30868|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001100;
  assign _0774_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30867|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001011;
  assign _0775_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30866|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001010;
  assign _0776_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30865|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001001;
  assign _0777_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30864|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10001000;
  assign _0778_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30863|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000111;
  assign _0779_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30862|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000110;
  assign _0780_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30861|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000101;
  assign _0781_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30860|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000100;
  assign _0782_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30859|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000011;
  assign _0783_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30858|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000010;
  assign _0784_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30857|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000001;
  assign _0785_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30856|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 8'b10000000;
  assign _0786_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30855|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111111;
  assign _0787_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30854|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111110;
  assign _0788_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30853|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111101;
  assign _0789_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30852|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111100;
  assign _0790_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30851|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111011;
  assign _0791_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30850|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111010;
  assign _0792_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30849|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111001;
  assign _0793_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30848|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1111000;
  assign _0794_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30847|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110111;
  assign _0795_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30846|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110110;
  assign _0796_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30845|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110101;
  assign _0797_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30844|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110100;
  assign _0798_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30843|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110011;
  assign _0799_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30842|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110010;
  assign _0800_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30841|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110001;
  assign _0801_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30840|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1110000;
  assign _0802_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30839|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101111;
  assign _0803_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30838|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101110;
  assign _0804_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30837|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101101;
  assign _0805_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30836|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101100;
  assign _0806_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30835|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101011;
  assign _0807_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30834|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101010;
  assign _0808_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30833|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101001;
  assign _0809_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30832|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1101000;
  assign _0810_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30831|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100111;
  assign _0811_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30830|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100110;
  assign _0812_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30829|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100101;
  assign _0813_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30828|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100100;
  assign _0814_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30827|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100011;
  assign _0815_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30826|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100010;
  assign _0816_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30825|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100001;
  assign _0817_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30824|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1100000;
  assign _0818_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30823|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011111;
  assign _0819_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30822|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011110;
  assign _0820_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30821|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011101;
  assign _0821_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30820|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011100;
  assign _0822_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30819|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011011;
  assign _0823_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30818|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011010;
  assign _0824_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30817|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011001;
  assign _0825_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30816|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1011000;
  assign _0826_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30815|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010111;
  assign _0827_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30814|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010110;
  assign _0828_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30813|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010101;
  assign _0829_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30812|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010100;
  assign _0830_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30811|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010011;
  assign _0831_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30810|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010010;
  assign _0832_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30809|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010001;
  assign _0833_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30808|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1010000;
  assign _0834_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30807|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001111;
  assign _0835_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30806|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001110;
  assign _0836_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30805|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001101;
  assign _0837_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30804|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001100;
  assign _0838_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30803|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001011;
  assign _0839_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30802|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001010;
  assign _0840_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30801|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001001;
  assign _0841_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30800|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1001000;
  assign _0842_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30799|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000111;
  assign _0843_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30798|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000110;
  assign _0844_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30797|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000101;
  assign _0845_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30796|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000100;
  assign _0846_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30795|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000011;
  assign _0847_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30794|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000010;
  assign _0848_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30793|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000001;
  assign _0849_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30792|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 7'b1000000;
  assign _0850_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30791|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111111;
  assign _0851_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30790|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111110;
  assign _0852_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30789|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111101;
  assign _0853_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30788|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111100;
  assign _0854_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30787|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111011;
  assign _0855_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30786|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111010;
  assign _0856_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30785|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111001;
  assign _0857_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30784|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b111000;
  assign _0858_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30783|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110111;
  assign _0859_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30782|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110110;
  assign _0860_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30781|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110101;
  assign _0861_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30780|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110100;
  assign _0862_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30779|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110011;
  assign _0863_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30778|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110010;
  assign _0864_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30777|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110001;
  assign _0865_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30776|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b110000;
  assign _0866_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30775|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101111;
  assign _0867_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30774|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101110;
  assign _0868_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30773|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101101;
  assign _0869_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30772|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101100;
  assign _0870_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30771|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101011;
  assign _0871_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30770|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101010;
  assign _0872_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30769|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101001;
  assign _0873_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30768|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b101000;
  assign _0874_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30767|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100111;
  assign _0875_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30766|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100110;
  assign _0876_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30765|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100101;
  assign _0877_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30764|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100100;
  assign _0878_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30763|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100011;
  assign _0879_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30762|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100010;
  assign _0880_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30761|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100001;
  assign _0881_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30760|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 6'b100000;
  assign _0882_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30759|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11111;
  assign _0883_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30758|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11110;
  assign _0884_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30757|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11101;
  assign _0885_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30756|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11100;
  assign _0886_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30755|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11011;
  assign _0887_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30754|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11010;
  assign _0888_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30753|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11001;
  assign _0889_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30752|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b11000;
  assign _0890_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30751|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10111;
  assign _0891_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30750|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10110;
  assign _0892_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30749|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10101;
  assign _0893_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30748|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10100;
  assign _0894_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30747|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10011;
  assign _0895_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30746|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10010;
  assign _0896_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30745|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10001;
  assign _0897_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30744|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 5'b10000;
  assign _0898_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30743|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1111;
  assign _0899_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30742|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1110;
  assign _0900_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30741|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1101;
  assign _0901_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30740|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1100;
  assign _0902_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30739|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1011;
  assign _0903_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30738|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1010;
  assign _0904_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30737|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1001;
  assign _0905_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30736|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 4'b1000;
  assign _0906_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30735|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 3'b111;
  assign _0907_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30734|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 3'b110;
  assign _0908_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30733|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 3'b101;
  assign _0909_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30732|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 3'b100;
  assign _0910_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30731|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 2'b11;
  assign _0911_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30730|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 2'b10;
  assign _0912_ = lut_in_addr3_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30729|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30728" *) 1'b1;
  function [15:0] _4003_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30461|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4003_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4003_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4003_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4003_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4003_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4003_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4003_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4003_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4003_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4003_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4003_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4003_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4003_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4003_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4003_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4003_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4003_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4003_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4003_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4003_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4003_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4003_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4003_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4003_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4003_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4003_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4003_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4003_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4003_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4003_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4003_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4003_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4003_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4003_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4003_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4003_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4003_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4003_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4003_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4003_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4003_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4003_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4003_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4003_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4003_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4003_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4003_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4003_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4003_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4003_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4003_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4003_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4003_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4003_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4003_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4003_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4003_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4003_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4003_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4003_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4003_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4003_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4003_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4003_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4003_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4003_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4003_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4003_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4003_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4003_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4003_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4003_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4003_ = b[4095:4080];
      default:
        _4003_ = a;
    endcase
  endfunction
  assign lo_data1_2 = _4003_(16'b0000000000000000, { REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_, _1032_, _1031_, _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0944_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_ });
  assign _0913_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30461|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 9'b100000000;
  assign _0914_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30460|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111111;
  assign _0915_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111110;
  assign _0916_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30458|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111101;
  assign _0917_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30457|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111100;
  assign _0918_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111011;
  assign _0919_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30455|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111010;
  assign _0920_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30454|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111001;
  assign _0921_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30453|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11111000;
  assign _0922_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30452|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110111;
  assign _0923_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30451|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110110;
  assign _0924_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30450|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110101;
  assign _0925_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30449|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110100;
  assign _0926_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30448|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110011;
  assign _0927_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110010;
  assign _0928_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30446|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110001;
  assign _0929_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30445|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11110000;
  assign _0930_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30444|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101111;
  assign _0931_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30443|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101110;
  assign _0932_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30442|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101101;
  assign _0933_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30441|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101100;
  assign _0934_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30440|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101011;
  assign _0935_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101010;
  assign _0936_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30438|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101001;
  assign _0937_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30437|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11101000;
  assign _0938_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30436|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100111;
  assign _0939_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30435|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100110;
  assign _0940_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30434|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100101;
  assign _0941_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30433|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100100;
  assign _0942_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30432|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100011;
  assign _0943_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30431|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100010;
  assign _0944_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30430|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100001;
  assign _0945_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30429|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11100000;
  assign _0946_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30428|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011111;
  assign _0947_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30427|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011110;
  assign _0948_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30426|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011101;
  assign _0949_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30425|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011100;
  assign _0950_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30424|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011011;
  assign _0951_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30423|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011010;
  assign _0952_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30422|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011001;
  assign _0953_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30421|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11011000;
  assign _0954_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30420|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010111;
  assign _0955_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30419|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010110;
  assign _0956_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30418|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010101;
  assign _0957_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30417|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010100;
  assign _0958_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30416|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010011;
  assign _0959_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30415|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010010;
  assign _0960_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30414|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010001;
  assign _0961_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30413|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11010000;
  assign _0962_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30412|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001111;
  assign _0963_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30411|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001110;
  assign _0964_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30410|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001101;
  assign _0965_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30409|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001100;
  assign _0966_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30408|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001011;
  assign _0967_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30407|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001010;
  assign _0968_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30406|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001001;
  assign _0969_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30405|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11001000;
  assign _0970_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30404|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000111;
  assign _0971_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30403|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000110;
  assign _0972_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30402|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000101;
  assign _0973_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30401|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000100;
  assign _0974_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30400|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000011;
  assign _0975_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30399|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000010;
  assign _0976_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30398|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000001;
  assign _0977_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30397|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b11000000;
  assign _0978_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30396|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111111;
  assign _0979_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30395|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111110;
  assign _0980_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30394|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111101;
  assign _0981_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30393|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111100;
  assign _0982_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30392|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111011;
  assign _0983_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30391|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111010;
  assign _0984_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30390|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111001;
  assign _0985_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30389|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10111000;
  assign _0986_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30388|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110111;
  assign _0987_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30387|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110110;
  assign _0988_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30386|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110101;
  assign _0989_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30385|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110100;
  assign _0990_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30384|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110011;
  assign _0991_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30383|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110010;
  assign _0992_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30382|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110001;
  assign _0993_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30381|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10110000;
  assign _0994_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30380|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101111;
  assign _0995_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30379|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101110;
  assign _0996_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30378|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101101;
  assign _0997_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30377|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101100;
  assign _0998_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30376|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101011;
  assign _0999_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30375|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101010;
  assign _1000_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30374|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101001;
  assign _1001_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30373|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10101000;
  assign _1002_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30372|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100111;
  assign _1003_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30371|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100110;
  assign _1004_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30370|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100101;
  assign _1005_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30369|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100100;
  assign _1006_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30368|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100011;
  assign _1007_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30367|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100010;
  assign _1008_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30366|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100001;
  assign _1009_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30365|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10100000;
  assign _1010_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30364|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011111;
  assign _1011_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30363|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011110;
  assign _1012_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30362|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011101;
  assign _1013_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30361|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011100;
  assign _1014_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30360|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011011;
  assign _1015_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30359|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011010;
  assign _1016_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30358|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011001;
  assign _1017_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30357|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10011000;
  assign _1018_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30356|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010111;
  assign _1019_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30355|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010110;
  assign _1020_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30354|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010101;
  assign _1021_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30353|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010100;
  assign _1022_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30352|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010011;
  assign _1023_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30351|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010010;
  assign _1024_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30350|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010001;
  assign _1025_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30349|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10010000;
  assign _1026_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30348|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001111;
  assign _1027_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30347|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001110;
  assign _1028_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30346|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001101;
  assign _1029_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30345|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001100;
  assign _1030_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30344|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001011;
  assign _1031_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30343|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001010;
  assign _1032_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30342|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001001;
  assign _1033_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30341|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10001000;
  assign _1034_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30340|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000111;
  assign _1035_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30339|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000110;
  assign _1036_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30338|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000101;
  assign _1037_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30337|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000100;
  assign _1038_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30336|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000011;
  assign _1039_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30335|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000010;
  assign _1040_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30334|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000001;
  assign _1041_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30333|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 8'b10000000;
  assign _1042_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30332|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111111;
  assign _1043_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30331|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111110;
  assign _1044_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30330|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111101;
  assign _1045_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30329|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111100;
  assign _1046_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30328|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111011;
  assign _1047_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30327|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111010;
  assign _1048_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30326|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111001;
  assign _1049_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30325|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1111000;
  assign _1050_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30324|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110111;
  assign _1051_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30323|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110110;
  assign _1052_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30322|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110101;
  assign _1053_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30321|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110100;
  assign _1054_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30320|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110011;
  assign _1055_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30319|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110010;
  assign _1056_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30318|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110001;
  assign _1057_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30317|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1110000;
  assign _1058_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30316|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101111;
  assign _1059_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30315|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101110;
  assign _1060_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30314|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101101;
  assign _1061_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30313|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101100;
  assign _1062_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30312|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101011;
  assign _1063_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30311|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101010;
  assign _1064_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30310|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101001;
  assign _1065_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30309|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1101000;
  assign _1066_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30308|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100111;
  assign _1067_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30307|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100110;
  assign _1068_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30306|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100101;
  assign _1069_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30305|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100100;
  assign _1070_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30304|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100011;
  assign _1071_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30303|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100010;
  assign _1072_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30302|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100001;
  assign _1073_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30301|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1100000;
  assign _1074_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30300|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011111;
  assign _1075_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30299|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011110;
  assign _1076_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30298|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011101;
  assign _1077_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30297|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011100;
  assign _1078_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30296|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011011;
  assign _1079_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30295|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011010;
  assign _1080_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30294|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011001;
  assign _1081_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30293|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1011000;
  assign _1082_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30292|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010111;
  assign _1083_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30291|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010110;
  assign _1084_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30290|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010101;
  assign _1085_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30289|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010100;
  assign _1086_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30288|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010011;
  assign _1087_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30287|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010010;
  assign _1088_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30286|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010001;
  assign _1089_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30285|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1010000;
  assign _1090_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30284|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001111;
  assign _1091_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30283|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001110;
  assign _1092_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30282|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001101;
  assign _1093_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30281|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001100;
  assign _1094_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30280|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001011;
  assign _1095_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30279|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001010;
  assign _1096_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30278|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001001;
  assign _1097_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30277|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1001000;
  assign _1098_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30276|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000111;
  assign _1099_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30275|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000110;
  assign _1100_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30274|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000101;
  assign _1101_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30273|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000100;
  assign _1102_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30272|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000011;
  assign _1103_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30271|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000010;
  assign _1104_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30270|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000001;
  assign _1105_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30269|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 7'b1000000;
  assign _1106_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30268|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111111;
  assign _1107_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30267|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111110;
  assign _1108_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30266|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111101;
  assign _1109_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30265|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111100;
  assign _1110_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30264|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111011;
  assign _1111_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30263|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111010;
  assign _1112_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30262|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111001;
  assign _1113_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30261|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b111000;
  assign _1114_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30260|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110111;
  assign _1115_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30259|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110110;
  assign _1116_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30258|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110101;
  assign _1117_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30257|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110100;
  assign _1118_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30256|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110011;
  assign _1119_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30255|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110010;
  assign _1120_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30254|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110001;
  assign _1121_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30253|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b110000;
  assign _1122_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30252|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101111;
  assign _1123_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30251|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101110;
  assign _1124_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30250|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101101;
  assign _1125_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30249|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101100;
  assign _1126_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30248|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101011;
  assign _1127_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30247|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101010;
  assign _1128_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30246|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101001;
  assign _1129_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30245|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b101000;
  assign _1130_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30244|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100111;
  assign _1131_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30243|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100110;
  assign _1132_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30242|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100101;
  assign _1133_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30241|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100100;
  assign _1134_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30240|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100011;
  assign _1135_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30239|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100010;
  assign _1136_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30238|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100001;
  assign _1137_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30237|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 6'b100000;
  assign _1138_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30236|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11111;
  assign _1139_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30235|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11110;
  assign _1140_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30234|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11101;
  assign _1141_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30233|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11100;
  assign _1142_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30232|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11011;
  assign _1143_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30231|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11010;
  assign _1144_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30230|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11001;
  assign _1145_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30229|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b11000;
  assign _1146_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30228|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10111;
  assign _1147_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30227|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10110;
  assign _1148_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30226|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10101;
  assign _1149_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30225|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10100;
  assign _1150_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30224|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10011;
  assign _1151_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30223|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10010;
  assign _1152_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30222|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10001;
  assign _1153_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30221|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 5'b10000;
  assign _1154_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30220|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1111;
  assign _1155_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30219|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1110;
  assign _1156_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30218|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1101;
  assign _1157_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30217|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1100;
  assign _1158_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30216|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1011;
  assign _1159_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30215|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1010;
  assign _1160_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30214|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1001;
  assign _1161_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30213|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 4'b1000;
  assign _1162_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30212|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 3'b111;
  assign _1163_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30211|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 3'b110;
  assign _1164_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30210|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 3'b101;
  assign _1165_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30209|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 3'b100;
  assign _1166_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30208|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 2'b11;
  assign _1167_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30207|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 2'b10;
  assign _1168_ = lut_in_addr2_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30206|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30205" *) 1'b1;
  function [15:0] _4260_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29938|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4260_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4260_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4260_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4260_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4260_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4260_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4260_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4260_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4260_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4260_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4260_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4260_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4260_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4260_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4260_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4260_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4260_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4260_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4260_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4260_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4260_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4260_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4260_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4260_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4260_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4260_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4260_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4260_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4260_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4260_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4260_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4260_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4260_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4260_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4260_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4260_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4260_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4260_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4260_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4260_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4260_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4260_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4260_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4260_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4260_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4260_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4260_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4260_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4260_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4260_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4260_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4260_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4260_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4260_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4260_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4260_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4260_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4260_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4260_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4260_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4260_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4260_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4260_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4260_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4260_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4260_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4260_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4260_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4260_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4260_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4260_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4260_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4260_ = b[4095:4080];
      default:
        _4260_ = a;
    endcase
  endfunction
  assign lo_data1_1 = _4260_(16'b0000000000000000, { REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_, _1290_, _1289_, _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_ });
  assign _1169_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29938|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 9'b100000000;
  assign _1170_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29937|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111111;
  assign _1171_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29936|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111110;
  assign _1172_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29935|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111101;
  assign _1173_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29934|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111100;
  assign _1174_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29933|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111011;
  assign _1175_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29932|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111010;
  assign _1176_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29931|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111001;
  assign _1177_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29930|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11111000;
  assign _1178_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29929|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110111;
  assign _1179_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29928|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110110;
  assign _1180_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29927|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110101;
  assign _1181_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29926|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110100;
  assign _1182_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29925|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110011;
  assign _1183_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29924|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110010;
  assign _1184_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29923|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110001;
  assign _1185_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29922|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11110000;
  assign _1186_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29921|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101111;
  assign _1187_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29920|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101110;
  assign _1188_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29919|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101101;
  assign _1189_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29918|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101100;
  assign _1190_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29917|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101011;
  assign _1191_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29916|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101010;
  assign _1192_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29915|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101001;
  assign _1193_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29914|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11101000;
  assign _1194_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29913|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100111;
  assign _1195_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29912|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100110;
  assign _1196_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29911|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100101;
  assign _1197_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29910|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100100;
  assign _1198_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29909|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100011;
  assign _1199_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29908|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100010;
  assign _1200_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29907|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100001;
  assign _1201_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29906|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11100000;
  assign _1202_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29905|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011111;
  assign _1203_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29904|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011110;
  assign _1204_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29903|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011101;
  assign _1205_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29902|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011100;
  assign _1206_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29901|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011011;
  assign _1207_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29900|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011010;
  assign _1208_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29899|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011001;
  assign _1209_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29898|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11011000;
  assign _1210_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29897|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010111;
  assign _1211_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29896|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010110;
  assign _1212_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29895|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010101;
  assign _1213_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29894|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010100;
  assign _1214_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29893|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010011;
  assign _1215_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29892|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010010;
  assign _1216_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29891|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010001;
  assign _1217_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29890|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11010000;
  assign _1218_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29889|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001111;
  assign _1219_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29888|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001110;
  assign _1220_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29887|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001101;
  assign _1221_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29886|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001100;
  assign _1222_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29885|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001011;
  assign _1223_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29884|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001010;
  assign _1224_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29883|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001001;
  assign _1225_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29882|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11001000;
  assign _1226_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29881|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000111;
  assign _1227_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29880|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000110;
  assign _1228_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29879|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000101;
  assign _1229_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29878|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000100;
  assign _1230_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29877|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000011;
  assign _1231_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29876|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000010;
  assign _1232_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29875|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000001;
  assign _1233_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29874|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b11000000;
  assign _1234_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29873|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111111;
  assign _1235_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29872|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111110;
  assign _1236_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29871|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111101;
  assign _1237_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29870|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111100;
  assign _1238_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29869|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111011;
  assign _1239_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29868|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111010;
  assign _1240_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29867|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111001;
  assign _1241_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29866|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10111000;
  assign _1242_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29865|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110111;
  assign _1243_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29864|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110110;
  assign _1244_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29863|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110101;
  assign _1245_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29862|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110100;
  assign _1246_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29861|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110011;
  assign _1247_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29860|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110010;
  assign _1248_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29859|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110001;
  assign _1249_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29858|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10110000;
  assign _1250_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29857|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101111;
  assign _1251_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29856|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101110;
  assign _1252_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29855|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101101;
  assign _1253_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29854|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101100;
  assign _1254_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29853|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101011;
  assign _1255_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29852|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101010;
  assign _1256_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29851|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101001;
  assign _1257_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29850|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10101000;
  assign _1258_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29849|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100111;
  assign _1259_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29848|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100110;
  assign _1260_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29847|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100101;
  assign _1261_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29846|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100100;
  assign _1262_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29845|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100011;
  assign _1263_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29844|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100010;
  assign _1264_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29843|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100001;
  assign _1265_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29842|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10100000;
  assign _1266_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29841|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011111;
  assign _1267_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29840|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011110;
  assign _1268_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29839|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011101;
  assign _1269_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29838|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011100;
  assign _1270_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29837|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011011;
  assign _1271_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29836|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011010;
  assign _1272_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29835|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011001;
  assign _1273_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29834|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10011000;
  assign _1274_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29833|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010111;
  assign _1275_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29832|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010110;
  assign _1276_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29831|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010101;
  assign _1277_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29830|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010100;
  assign _1278_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29829|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010011;
  assign _1279_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29828|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010010;
  assign _1280_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29827|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010001;
  assign _1281_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29826|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10010000;
  assign _1282_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29825|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001111;
  assign _1283_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29824|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001110;
  assign _1284_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29823|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001101;
  assign _1285_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29822|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001100;
  assign _1286_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29821|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001011;
  assign _1287_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29820|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001010;
  assign _1288_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29819|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001001;
  assign _1289_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29818|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10001000;
  assign _1290_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29817|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000111;
  assign _1291_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29816|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000110;
  assign _1292_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29815|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000101;
  assign _1293_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29814|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000100;
  assign _1294_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29813|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000011;
  assign _1295_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29812|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000010;
  assign _1296_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29811|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000001;
  assign _1297_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29810|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 8'b10000000;
  assign _1298_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29809|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111111;
  assign _1299_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29808|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111110;
  assign _1300_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29807|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111101;
  assign _1301_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29806|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111100;
  assign _1302_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29805|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111011;
  assign _1303_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29804|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111010;
  assign _1304_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29803|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111001;
  assign _1305_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29802|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1111000;
  assign _1306_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29801|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110111;
  assign _1307_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29800|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110110;
  assign _1308_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29799|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110101;
  assign _1309_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29798|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110100;
  assign _1310_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29797|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110011;
  assign _1311_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29796|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110010;
  assign _1312_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29795|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110001;
  assign _1313_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29794|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1110000;
  assign _1314_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29793|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101111;
  assign _1315_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29792|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101110;
  assign _1316_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29791|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101101;
  assign _1317_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29790|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101100;
  assign _1318_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29789|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101011;
  assign _1319_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29788|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101010;
  assign _1320_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29787|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101001;
  assign _1321_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29786|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1101000;
  assign _1322_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29785|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100111;
  assign _1323_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29784|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100110;
  assign _1324_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29783|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100101;
  assign _1325_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29782|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100100;
  assign _1326_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29781|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100011;
  assign _1327_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29780|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100010;
  assign _1328_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29779|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100001;
  assign _1329_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29778|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1100000;
  assign _1330_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29777|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011111;
  assign _1331_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29776|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011110;
  assign _1332_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29775|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011101;
  assign _1333_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29774|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011100;
  assign _1334_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29773|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011011;
  assign _1335_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29772|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011010;
  assign _1336_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29771|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011001;
  assign _1337_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29770|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1011000;
  assign _1338_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29769|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010111;
  assign _1339_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29768|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010110;
  assign _1340_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29767|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010101;
  assign _1341_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29766|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010100;
  assign _1342_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29765|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010011;
  assign _1343_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29764|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010010;
  assign _1344_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29763|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010001;
  assign _1345_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29762|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1010000;
  assign _1346_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29761|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001111;
  assign _1347_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29760|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001110;
  assign _1348_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29759|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001101;
  assign _1349_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29758|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001100;
  assign _1350_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29757|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001011;
  assign _1351_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29756|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001010;
  assign _1352_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29755|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001001;
  assign _1353_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29754|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1001000;
  assign _1354_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29753|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000111;
  assign _1355_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29752|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000110;
  assign _1356_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29751|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000101;
  assign _1357_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29750|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000100;
  assign _1358_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29749|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000011;
  assign _1359_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29748|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000010;
  assign _1360_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29747|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000001;
  assign _1361_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29746|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 7'b1000000;
  assign _1362_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29745|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111111;
  assign _1363_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29744|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111110;
  assign _1364_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29743|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111101;
  assign _1365_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29742|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111100;
  assign _1366_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29741|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111011;
  assign _1367_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29740|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111010;
  assign _1368_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29739|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111001;
  assign _1369_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29738|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b111000;
  assign _1370_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29737|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110111;
  assign _1371_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29736|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110110;
  assign _1372_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29735|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110101;
  assign _1373_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29734|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110100;
  assign _1374_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29733|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110011;
  assign _1375_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29732|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110010;
  assign _1376_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29731|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110001;
  assign _1377_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29730|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b110000;
  assign _1378_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29729|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101111;
  assign _1379_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29728|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101110;
  assign _1380_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29727|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101101;
  assign _1381_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29726|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101100;
  assign _1382_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29725|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101011;
  assign _1383_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29724|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101010;
  assign _1384_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29723|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101001;
  assign _1385_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29722|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b101000;
  assign _1386_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29721|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100111;
  assign _1387_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29720|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100110;
  assign _1388_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29719|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100101;
  assign _1389_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29718|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100100;
  assign _1390_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29717|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100011;
  assign _1391_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29716|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100010;
  assign _1392_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29715|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100001;
  assign _1393_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29714|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 6'b100000;
  assign _1394_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29713|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11111;
  assign _1395_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29712|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11110;
  assign _1396_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29711|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11101;
  assign _1397_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29710|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11100;
  assign _1398_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29709|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11011;
  assign _1399_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29708|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11010;
  assign _1400_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29707|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11001;
  assign _1401_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29706|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b11000;
  assign _1402_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29705|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10111;
  assign _1403_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29704|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10110;
  assign _1404_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29703|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10101;
  assign _1405_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29702|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10100;
  assign _1406_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29701|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10011;
  assign _1407_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29700|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10010;
  assign _1408_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29699|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10001;
  assign _1409_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29698|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 5'b10000;
  assign _1410_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29697|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1111;
  assign _1411_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29696|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1110;
  assign _1412_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29695|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1101;
  assign _1413_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29694|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1100;
  assign _1414_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29693|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1011;
  assign _1415_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29692|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1010;
  assign _1416_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29691|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1001;
  assign _1417_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29690|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 4'b1000;
  assign _1418_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29689|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 3'b111;
  assign _1419_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29688|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 3'b110;
  assign _1420_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29687|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 3'b101;
  assign _1421_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29686|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 3'b100;
  assign _1422_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29685|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 2'b11;
  assign _1423_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29684|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 2'b10;
  assign _1424_ = lut_in_addr1_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29683|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29682" *) 1'b1;
  function [15:0] _4517_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29415|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4517_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4517_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4517_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4517_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4517_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4517_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4517_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4517_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4517_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4517_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4517_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4517_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4517_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4517_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4517_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4517_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4517_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4517_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4517_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4517_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4517_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4517_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4517_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4517_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4517_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4517_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4517_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4517_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4517_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4517_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4517_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4517_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4517_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4517_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4517_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4517_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4517_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4517_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4517_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4517_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4517_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4517_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4517_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4517_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4517_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4517_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4517_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4517_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4517_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4517_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4517_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4517_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4517_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4517_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4517_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4517_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4517_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4517_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4517_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4517_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4517_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4517_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4517_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4517_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4517_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4517_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4517_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4517_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4517_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4517_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4517_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4517_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4517_ = b[4095:4080];
      default:
        _4517_ = a;
    endcase
  endfunction
  assign lo_data1_0 = _4517_(16'b0000000000000000, { REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_, _1548_, _1547_, _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_, _1470_, _1469_, _1468_, _1467_, _1466_, _1465_, _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_ });
  assign _1425_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29415|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 9'b100000000;
  assign _1426_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29414|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111111;
  assign _1427_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29413|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111110;
  assign _1428_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29412|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111101;
  assign _1429_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29411|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111100;
  assign _1430_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29410|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111011;
  assign _1431_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29409|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111010;
  assign _1432_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29408|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111001;
  assign _1433_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29407|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11111000;
  assign _1434_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29406|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110111;
  assign _1435_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29405|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110110;
  assign _1436_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29404|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110101;
  assign _1437_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29403|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110100;
  assign _1438_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29402|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110011;
  assign _1439_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29401|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110010;
  assign _1440_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29400|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110001;
  assign _1441_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29399|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11110000;
  assign _1442_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29398|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101111;
  assign _1443_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29397|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101110;
  assign _1444_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29396|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101101;
  assign _1445_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29395|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101100;
  assign _1446_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29394|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101011;
  assign _1447_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29393|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101010;
  assign _1448_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29392|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101001;
  assign _1449_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29391|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11101000;
  assign _1450_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29390|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100111;
  assign _1451_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29389|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100110;
  assign _1452_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29388|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100101;
  assign _1453_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29387|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100100;
  assign _1454_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29386|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100011;
  assign _1455_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29385|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100010;
  assign _1456_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29384|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100001;
  assign _1457_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29383|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11100000;
  assign _1458_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29382|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011111;
  assign _1459_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29381|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011110;
  assign _1460_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29380|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011101;
  assign _1461_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29379|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011100;
  assign _1462_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29378|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011011;
  assign _1463_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29377|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011010;
  assign _1464_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29376|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011001;
  assign _1465_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29375|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11011000;
  assign _1466_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29374|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010111;
  assign _1467_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29373|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010110;
  assign _1468_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29372|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010101;
  assign _1469_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29371|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010100;
  assign _1470_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29370|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010011;
  assign _1471_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29369|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010010;
  assign _1472_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29368|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010001;
  assign _1473_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29367|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11010000;
  assign _1474_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29366|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001111;
  assign _1475_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29365|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001110;
  assign _1476_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29364|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001101;
  assign _1477_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29363|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001100;
  assign _1478_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29362|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001011;
  assign _1479_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29361|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001010;
  assign _1480_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29360|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001001;
  assign _1481_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29359|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11001000;
  assign _1482_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29358|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000111;
  assign _1483_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29357|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000110;
  assign _1484_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29356|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000101;
  assign _1485_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29355|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000100;
  assign _1486_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29354|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000011;
  assign _1487_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29353|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000010;
  assign _1488_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29352|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000001;
  assign _1489_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29351|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b11000000;
  assign _1490_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29350|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111111;
  assign _1491_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29349|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111110;
  assign _1492_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29348|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111101;
  assign _1493_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29347|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111100;
  assign _1494_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29346|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111011;
  assign _1495_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29345|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111010;
  assign _1496_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29344|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111001;
  assign _1497_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29343|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10111000;
  assign _1498_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29342|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110111;
  assign _1499_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29341|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110110;
  assign _1500_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29340|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110101;
  assign _1501_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29339|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110100;
  assign _1502_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29338|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110011;
  assign _1503_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29337|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110010;
  assign _1504_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29336|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110001;
  assign _1505_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29335|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10110000;
  assign _1506_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29334|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101111;
  assign _1507_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29333|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101110;
  assign _1508_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29332|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101101;
  assign _1509_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29331|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101100;
  assign _1510_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29330|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101011;
  assign _1511_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29329|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101010;
  assign _1512_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29328|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101001;
  assign _1513_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29327|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10101000;
  assign _1514_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29326|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100111;
  assign _1515_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29325|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100110;
  assign _1516_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29324|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100101;
  assign _1517_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29323|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100100;
  assign _1518_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29322|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100011;
  assign _1519_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29321|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100010;
  assign _1520_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29320|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100001;
  assign _1521_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29319|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10100000;
  assign _1522_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29318|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011111;
  assign _1523_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29317|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011110;
  assign _1524_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29316|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011101;
  assign _1525_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29315|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011100;
  assign _1526_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29314|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011011;
  assign _1527_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29313|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011010;
  assign _1528_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29312|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011001;
  assign _1529_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29311|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10011000;
  assign _1530_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29310|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010111;
  assign _1531_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29309|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010110;
  assign _1532_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29308|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010101;
  assign _1533_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29307|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010100;
  assign _1534_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29306|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010011;
  assign _1535_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29305|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010010;
  assign _1536_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29304|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010001;
  assign _1537_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29303|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10010000;
  assign _1538_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29302|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001111;
  assign _1539_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29301|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001110;
  assign _1540_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29300|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001101;
  assign _1541_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29299|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001100;
  assign _1542_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29298|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001011;
  assign _1543_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29297|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001010;
  assign _1544_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29296|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001001;
  assign _1545_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29295|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10001000;
  assign _1546_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29294|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000111;
  assign _1547_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29293|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000110;
  assign _1548_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29292|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000101;
  assign _1549_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29291|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000100;
  assign _1550_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29290|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000011;
  assign _1551_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29289|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000010;
  assign _1552_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29288|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000001;
  assign _1553_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29287|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 8'b10000000;
  assign _1554_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29286|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111111;
  assign _1555_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29285|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111110;
  assign _1556_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29284|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111101;
  assign _1557_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29283|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111100;
  assign _1558_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29282|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111011;
  assign _1559_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29281|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111010;
  assign _1560_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29280|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111001;
  assign _1561_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29279|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1111000;
  assign _1562_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29278|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110111;
  assign _1563_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29277|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110110;
  assign _1564_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29276|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110101;
  assign _1565_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29275|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110100;
  assign _1566_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29274|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110011;
  assign _1567_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29273|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110010;
  assign _1568_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29272|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110001;
  assign _1569_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29271|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1110000;
  assign _1570_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29270|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101111;
  assign _1571_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29269|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101110;
  assign _1572_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29268|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101101;
  assign _1573_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29267|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101100;
  assign _1574_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29266|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101011;
  assign _1575_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29265|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101010;
  assign _1576_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29264|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101001;
  assign _1577_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29263|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1101000;
  assign _1578_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29262|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100111;
  assign _1579_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29261|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100110;
  assign _1580_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29260|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100101;
  assign _1581_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29259|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100100;
  assign _1582_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29258|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100011;
  assign _1583_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29257|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100010;
  assign _1584_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29256|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100001;
  assign _1585_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29255|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1100000;
  assign _1586_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29254|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011111;
  assign _1587_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29253|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011110;
  assign _1588_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29252|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011101;
  assign _1589_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29251|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011100;
  assign _1590_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29250|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011011;
  assign _1591_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29249|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011010;
  assign _1592_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29248|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011001;
  assign _1593_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29247|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1011000;
  assign _1594_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29246|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010111;
  assign _1595_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29245|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010110;
  assign _1596_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29244|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010101;
  assign _1597_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29243|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010100;
  assign _1598_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29242|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010011;
  assign _1599_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29241|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010010;
  assign _1600_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29240|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010001;
  assign _1601_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29239|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1010000;
  assign _1602_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29238|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001111;
  assign _1603_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29237|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001110;
  assign _1604_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29236|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001101;
  assign _1605_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29235|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001100;
  assign _1606_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29234|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001011;
  assign _1607_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29233|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001010;
  assign _1608_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29232|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001001;
  assign _1609_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29231|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1001000;
  assign _1610_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29230|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000111;
  assign _1611_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29229|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000110;
  assign _1612_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29228|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000101;
  assign _1613_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29227|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000100;
  assign _1614_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29226|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000011;
  assign _1615_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29225|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000010;
  assign _1616_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29224|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000001;
  assign _1617_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29223|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 7'b1000000;
  assign _1618_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29222|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111111;
  assign _1619_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29221|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111110;
  assign _1620_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29220|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111101;
  assign _1621_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29219|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111100;
  assign _1622_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29218|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111011;
  assign _1623_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29217|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111010;
  assign _1624_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29216|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111001;
  assign _1625_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29215|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b111000;
  assign _1626_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29214|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110111;
  assign _1627_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29213|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110110;
  assign _1628_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29212|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110101;
  assign _1629_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29211|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110100;
  assign _1630_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29210|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110011;
  assign _1631_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29209|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110010;
  assign _1632_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29208|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110001;
  assign _1633_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29207|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b110000;
  assign _1634_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29206|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101111;
  assign _1635_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29205|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101110;
  assign _1636_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29204|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101101;
  assign _1637_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29203|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101100;
  assign _1638_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29202|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101011;
  assign _1639_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29201|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101010;
  assign _1640_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29200|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101001;
  assign _1641_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29199|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b101000;
  assign _1642_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29198|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100111;
  assign _1643_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29197|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100110;
  assign _1644_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29196|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100101;
  assign _1645_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29195|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100100;
  assign _1646_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29194|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100011;
  assign _1647_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29193|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100010;
  assign _1648_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29192|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100001;
  assign _1649_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29191|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 6'b100000;
  assign _1650_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29190|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11111;
  assign _1651_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29189|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11110;
  assign _1652_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29188|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11101;
  assign _1653_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29187|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11100;
  assign _1654_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29186|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11011;
  assign _1655_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29185|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11010;
  assign _1656_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29184|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11001;
  assign _1657_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29183|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b11000;
  assign _1658_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29182|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10111;
  assign _1659_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29181|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10110;
  assign _1660_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29180|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10101;
  assign _1661_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29179|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10100;
  assign _1662_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29178|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10011;
  assign _1663_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29177|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10010;
  assign _1664_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29176|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10001;
  assign _1665_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29175|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 5'b10000;
  assign _1666_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29174|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1111;
  assign _1667_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29173|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1110;
  assign _1668_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29172|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1101;
  assign _1669_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29171|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1100;
  assign _1670_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29170|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1011;
  assign _1671_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29169|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1010;
  assign _1672_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29168|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1001;
  assign _1673_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29167|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 4'b1000;
  assign _1674_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29166|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 3'b111;
  assign _1675_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29165|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 3'b110;
  assign _1676_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29164|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 3'b101;
  assign _1677_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29163|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 3'b100;
  assign _1678_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29162|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 2'b11;
  assign _1679_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29161|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 2'b10;
  assign _1680_ = lut_in_addr0_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29160|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:29159" *) 1'b1;
  function [15:0] _4774_;
    input [15:0] a;
    input [4111:0] b;
    input [256:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28892|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *)
    (* parallel_case *)
    casez (s)
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4774_ = b[15:0];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4774_ = b[31:16];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4774_ = b[47:32];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4774_ = b[63:48];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4774_ = b[79:64];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4774_ = b[95:80];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4774_ = b[111:96];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4774_ = b[127:112];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4774_ = b[143:128];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4774_ = b[159:144];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4774_ = b[175:160];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4774_ = b[191:176];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4774_ = b[207:192];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4774_ = b[223:208];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4774_ = b[239:224];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4774_ = b[255:240];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4774_ = b[271:256];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4774_ = b[287:272];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4774_ = b[303:288];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4774_ = b[319:304];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4774_ = b[335:320];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4774_ = b[351:336];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4774_ = b[367:352];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4774_ = b[383:368];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4774_ = b[399:384];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4774_ = b[415:400];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4774_ = b[431:416];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4774_ = b[447:432];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4774_ = b[463:448];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4774_ = b[479:464];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4774_ = b[495:480];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4774_ = b[511:496];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4774_ = b[527:512];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4774_ = b[543:528];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4774_ = b[559:544];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4774_ = b[575:560];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4774_ = b[591:576];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4774_ = b[607:592];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4774_ = b[623:608];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4774_ = b[639:624];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4774_ = b[655:640];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4774_ = b[671:656];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4774_ = b[687:672];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4774_ = b[703:688];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4774_ = b[719:704];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4774_ = b[735:720];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4774_ = b[751:736];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4774_ = b[767:752];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4774_ = b[783:768];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4774_ = b[799:784];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4774_ = b[815:800];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4774_ = b[831:816];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4774_ = b[847:832];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4774_ = b[863:848];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4774_ = b[879:864];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4774_ = b[895:880];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4774_ = b[911:896];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4774_ = b[927:912];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4774_ = b[943:928];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4774_ = b[959:944];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4774_ = b[975:960];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4774_ = b[991:976];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4774_ = b[1007:992];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4774_ = b[1023:1008];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4774_ = b[1039:1024];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4774_ = b[1055:1040];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4774_ = b[1071:1056];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4774_ = b[1087:1072];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4774_ = b[1103:1088];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4774_ = b[1119:1104];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4774_ = b[1135:1120];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4774_ = b[1151:1136];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1167:1152];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1183:1168];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1199:1184];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1215:1200];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1231:1216];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1247:1232];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1263:1248];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1279:1264];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1295:1280];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1311:1296];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1327:1312];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1343:1328];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1359:1344];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1375:1360];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1391:1376];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1407:1392];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1423:1408];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1439:1424];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1455:1440];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1471:1456];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1487:1472];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1503:1488];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1519:1504];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1535:1520];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1551:1536];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1567:1552];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1583:1568];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1599:1584];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1615:1600];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1631:1616];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1647:1632];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1663:1648];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1679:1664];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1695:1680];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1711:1696];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1727:1712];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1743:1728];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1759:1744];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1775:1760];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1791:1776];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1807:1792];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1823:1808];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1839:1824];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1855:1840];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1871:1856];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1887:1872];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1903:1888];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1919:1904];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1935:1920];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1951:1936];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1967:1952];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1983:1968];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[1999:1984];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2015:2000];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2031:2016];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2047:2032];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2063:2048];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2079:2064];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2095:2080];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2111:2096];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2127:2112];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2143:2128];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2159:2144];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2175:2160];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2191:2176];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2207:2192];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2223:2208];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2239:2224];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2255:2240];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2271:2256];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2287:2272];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2303:2288];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2319:2304];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2335:2320];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2351:2336];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2367:2352];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2383:2368];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2399:2384];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2415:2400];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2431:2416];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2447:2432];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2463:2448];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2479:2464];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2495:2480];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2511:2496];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2527:2512];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2543:2528];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2559:2544];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2575:2560];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2591:2576];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2607:2592];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2623:2608];
      257'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2639:2624];
      257'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2655:2640];
      257'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2671:2656];
      257'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2687:2672];
      257'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2703:2688];
      257'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2719:2704];
      257'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2735:2720];
      257'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2751:2736];
      257'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2767:2752];
      257'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2783:2768];
      257'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2799:2784];
      257'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2815:2800];
      257'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2831:2816];
      257'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2847:2832];
      257'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2863:2848];
      257'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2879:2864];
      257'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2895:2880];
      257'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2911:2896];
      257'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2927:2912];
      257'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2943:2928];
      257'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2959:2944];
      257'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2975:2960];
      257'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[2991:2976];
      257'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3007:2992];
      257'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3023:3008];
      257'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3039:3024];
      257'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3055:3040];
      257'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3071:3056];
      257'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3087:3072];
      257'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3103:3088];
      257'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3119:3104];
      257'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3135:3120];
      257'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3151:3136];
      257'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3167:3152];
      257'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3183:3168];
      257'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3199:3184];
      257'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3215:3200];
      257'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3231:3216];
      257'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3247:3232];
      257'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3263:3248];
      257'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3279:3264];
      257'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3295:3280];
      257'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3311:3296];
      257'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3327:3312];
      257'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3343:3328];
      257'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3359:3344];
      257'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3375:3360];
      257'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3391:3376];
      257'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3407:3392];
      257'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3423:3408];
      257'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3439:3424];
      257'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3455:3440];
      257'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3471:3456];
      257'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3487:3472];
      257'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3503:3488];
      257'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3519:3504];
      257'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3535:3520];
      257'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3551:3536];
      257'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3567:3552];
      257'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3583:3568];
      257'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3599:3584];
      257'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3615:3600];
      257'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3631:3616];
      257'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3647:3632];
      257'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3663:3648];
      257'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3679:3664];
      257'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3695:3680];
      257'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3711:3696];
      257'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3727:3712];
      257'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3743:3728];
      257'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3759:3744];
      257'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3775:3760];
      257'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3791:3776];
      257'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3807:3792];
      257'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3823:3808];
      257'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3839:3824];
      257'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3855:3840];
      257'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3871:3856];
      257'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3887:3872];
      257'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3903:3888];
      257'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3919:3904];
      257'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3935:3920];
      257'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3951:3936];
      257'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3967:3952];
      257'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3983:3968];
      257'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[3999:3984];
      257'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4015:4000];
      257'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4031:4016];
      257'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4047:4032];
      257'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4063:4048];
      257'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4079:4064];
      257'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4095:4080];
      257'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4774_ = b[4111:4096];
      default:
        _4774_ = a;
    endcase
  endfunction
  assign lo_data0_3 = _4774_(16'b0000000000000000, { REG_lo_0, REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_, _1806_, _1805_, _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_, _1733_, _1732_, _1731_, _1730_, _1729_, _1728_, _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_ });
  assign _1681_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28892|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 9'b100000000;
  assign _1682_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28891|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111111;
  assign _1683_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28890|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111110;
  assign _1684_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28889|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111101;
  assign _1685_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28888|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111100;
  assign _1686_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28887|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111011;
  assign _1687_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28886|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111010;
  assign _1688_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28885|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111001;
  assign _1689_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28884|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11111000;
  assign _1690_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28883|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110111;
  assign _1691_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28882|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110110;
  assign _1692_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28881|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110101;
  assign _1693_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28880|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110100;
  assign _1694_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28879|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110011;
  assign _1695_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28878|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110010;
  assign _1696_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28877|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110001;
  assign _1697_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28876|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11110000;
  assign _1698_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28875|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101111;
  assign _1699_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28874|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101110;
  assign _1700_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28873|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101101;
  assign _1701_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28872|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101100;
  assign _1702_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28871|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101011;
  assign _1703_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28870|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101010;
  assign _1704_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28869|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101001;
  assign _1705_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28868|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11101000;
  assign _1706_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28867|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100111;
  assign _1707_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28866|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100110;
  assign _1708_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28865|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100101;
  assign _1709_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28864|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100100;
  assign _1710_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28863|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100011;
  assign _1711_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28862|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100010;
  assign _1712_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28861|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100001;
  assign _1713_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28860|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11100000;
  assign _1714_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28859|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011111;
  assign _1715_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28858|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011110;
  assign _1716_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28857|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011101;
  assign _1717_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28856|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011100;
  assign _1718_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28855|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011011;
  assign _1719_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28854|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011010;
  assign _1720_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28853|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011001;
  assign _1721_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28852|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11011000;
  assign _1722_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28851|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010111;
  assign _1723_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28850|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010110;
  assign _1724_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28849|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010101;
  assign _1725_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28848|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010100;
  assign _1726_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28847|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010011;
  assign _1727_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28846|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010010;
  assign _1728_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28845|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010001;
  assign _1729_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28844|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11010000;
  assign _1730_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28843|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001111;
  assign _1731_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28842|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001110;
  assign _1732_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28841|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001101;
  assign _1733_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28840|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001100;
  assign _1734_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28839|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001011;
  assign _1735_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28838|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001010;
  assign _1736_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28837|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001001;
  assign _1737_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28836|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11001000;
  assign _1738_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28835|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000111;
  assign _1739_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28834|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000110;
  assign _1740_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28833|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000101;
  assign _1741_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28832|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000100;
  assign _1742_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28831|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000011;
  assign _1743_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28830|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000010;
  assign _1744_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28829|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000001;
  assign _1745_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28828|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b11000000;
  assign _1746_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28827|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111111;
  assign _1747_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28826|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111110;
  assign _1748_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28825|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111101;
  assign _1749_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28824|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111100;
  assign _1750_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28823|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111011;
  assign _1751_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28822|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111010;
  assign _1752_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28821|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111001;
  assign _1753_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28820|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10111000;
  assign _1754_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28819|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110111;
  assign _1755_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28818|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110110;
  assign _1756_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28817|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110101;
  assign _1757_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28816|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110100;
  assign _1758_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28815|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110011;
  assign _1759_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28814|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110010;
  assign _1760_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28813|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110001;
  assign _1761_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28812|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10110000;
  assign _1762_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28811|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101111;
  assign _1763_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28810|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101110;
  assign _1764_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28809|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101101;
  assign _1765_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28808|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101100;
  assign _1766_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28807|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101011;
  assign _1767_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28806|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101010;
  assign _1768_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28805|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101001;
  assign _1769_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28804|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10101000;
  assign _1770_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28803|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100111;
  assign _1771_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28802|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100110;
  assign _1772_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28801|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100101;
  assign _1773_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28800|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100100;
  assign _1774_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28799|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100011;
  assign _1775_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28798|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100010;
  assign _1776_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28797|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100001;
  assign _1777_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28796|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10100000;
  assign _1778_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28795|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011111;
  assign _1779_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28794|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011110;
  assign _1780_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28793|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011101;
  assign _1781_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28792|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011100;
  assign _1782_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28791|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011011;
  assign _1783_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28790|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011010;
  assign _1784_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28789|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011001;
  assign _1785_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28788|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10011000;
  assign _1786_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28787|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010111;
  assign _1787_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28786|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010110;
  assign _1788_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28785|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010101;
  assign _1789_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28784|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010100;
  assign _1790_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28783|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010011;
  assign _1791_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28782|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010010;
  assign _1792_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28781|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010001;
  assign _1793_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28780|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10010000;
  assign _1794_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28779|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001111;
  assign _1795_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28778|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001110;
  assign _1796_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28777|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001101;
  assign _1797_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28776|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001100;
  assign _1798_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28775|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001011;
  assign _1799_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28774|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001010;
  assign _1800_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28773|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001001;
  assign _1801_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28772|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10001000;
  assign _1802_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28771|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000111;
  assign _1803_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28770|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000110;
  assign _1804_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28769|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000101;
  assign _1805_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28768|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000100;
  assign _1806_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28767|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000011;
  assign _1807_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28766|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000010;
  assign _1808_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28765|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000001;
  assign _1809_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28764|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 8'b10000000;
  assign _1810_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28763|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111111;
  assign _1811_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28762|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111110;
  assign _1812_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28761|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111101;
  assign _1813_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28760|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111100;
  assign _1814_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28759|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111011;
  assign _1815_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28758|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111010;
  assign _1816_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28757|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111001;
  assign _1817_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28756|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1111000;
  assign _1818_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28755|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110111;
  assign _1819_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28754|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110110;
  assign _1820_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28753|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110101;
  assign _1821_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28752|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110100;
  assign _1822_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28751|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110011;
  assign _1823_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28750|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110010;
  assign _1824_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28749|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110001;
  assign _1825_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28748|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1110000;
  assign _1826_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28747|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101111;
  assign _1827_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28746|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101110;
  assign _1828_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28745|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101101;
  assign _1829_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28744|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101100;
  assign _1830_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28743|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101011;
  assign _1831_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28742|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101010;
  assign _1832_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28741|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101001;
  assign _1833_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28740|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1101000;
  assign _1834_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28739|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100111;
  assign _1835_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28738|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100110;
  assign _1836_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28737|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100101;
  assign _1837_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28736|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100100;
  assign _1838_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28735|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100011;
  assign _1839_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28734|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100010;
  assign _1840_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28733|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100001;
  assign _1841_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28732|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1100000;
  assign _1842_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28731|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011111;
  assign _1843_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28730|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011110;
  assign _1844_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28729|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011101;
  assign _1845_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28728|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011100;
  assign _1846_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28727|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011011;
  assign _1847_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28726|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011010;
  assign _1848_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28725|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011001;
  assign _1849_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28724|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1011000;
  assign _1850_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28723|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010111;
  assign _1851_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28722|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010110;
  assign _1852_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28721|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010101;
  assign _1853_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28720|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010100;
  assign _1854_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28719|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010011;
  assign _1855_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28718|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010010;
  assign _1856_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28717|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010001;
  assign _1857_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28716|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1010000;
  assign _1858_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28715|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001111;
  assign _1859_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28714|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001110;
  assign _1860_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28713|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001101;
  assign _1861_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28712|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001100;
  assign _1862_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28711|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001011;
  assign _1863_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28710|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001010;
  assign _1864_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28709|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001001;
  assign _1865_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28708|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1001000;
  assign _1866_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28707|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000111;
  assign _1867_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28706|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000110;
  assign _1868_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28705|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000101;
  assign _1869_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28704|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000100;
  assign _1870_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28703|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000011;
  assign _1871_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28702|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000010;
  assign _1872_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28701|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000001;
  assign _1873_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28700|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 7'b1000000;
  assign _1874_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28699|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111111;
  assign _1875_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28698|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111110;
  assign _1876_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28697|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111101;
  assign _1877_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28696|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111100;
  assign _1878_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28695|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111011;
  assign _1879_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28694|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111010;
  assign _1880_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28693|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111001;
  assign _1881_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28692|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b111000;
  assign _1882_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28691|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110111;
  assign _1883_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28690|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110110;
  assign _1884_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28689|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110101;
  assign _1885_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28688|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110100;
  assign _1886_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28687|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110011;
  assign _1887_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28686|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110010;
  assign _1888_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28685|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110001;
  assign _1889_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28684|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b110000;
  assign _1890_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28683|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101111;
  assign _1891_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28682|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101110;
  assign _1892_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28681|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101101;
  assign _1893_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28680|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101100;
  assign _1894_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28679|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101011;
  assign _1895_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28678|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101010;
  assign _1896_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28677|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101001;
  assign _1897_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28676|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b101000;
  assign _1898_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28675|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100111;
  assign _1899_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28674|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100110;
  assign _1900_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28673|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100101;
  assign _1901_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28672|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100100;
  assign _1902_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28671|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100011;
  assign _1903_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28670|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100010;
  assign _1904_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28669|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100001;
  assign _1905_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28668|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 6'b100000;
  assign _1906_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28667|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11111;
  assign _1907_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28666|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11110;
  assign _1908_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28665|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11101;
  assign _1909_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28664|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11100;
  assign _1910_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28663|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11011;
  assign _1911_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28662|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11010;
  assign _1912_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28661|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11001;
  assign _1913_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28660|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b11000;
  assign _1914_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10111;
  assign _1915_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28658|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10110;
  assign _1916_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28657|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10101;
  assign _1917_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28656|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10100;
  assign _1918_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28655|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10011;
  assign _1919_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28654|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10010;
  assign _1920_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28653|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10001;
  assign _1921_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28652|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 5'b10000;
  assign _1922_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28651|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1111;
  assign _1923_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28650|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1110;
  assign _1924_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28649|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1101;
  assign _1925_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28648|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1100;
  assign _1926_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28647|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1011;
  assign _1927_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28646|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1010;
  assign _1928_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28645|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1001;
  assign _1929_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28644|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 4'b1000;
  assign _1930_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28643|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 3'b111;
  assign _1931_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 3'b110;
  assign _1932_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28641|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 3'b101;
  assign _1933_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28640|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 3'b100;
  assign _1934_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28639|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 2'b11;
  assign _1935_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28638|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 2'b10;
  assign _1936_ = p1_pipe_data[315:307] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28637|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) 1'b1;
  assign _1937_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28636|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28635" *) p1_pipe_data[315:307];
  function [15:0] _5032_;
    input [15:0] a;
    input [4111:0] b;
    input [256:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28367|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *)
    (* parallel_case *)
    casez (s)
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5032_ = b[15:0];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5032_ = b[31:16];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5032_ = b[47:32];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5032_ = b[63:48];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5032_ = b[79:64];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5032_ = b[95:80];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5032_ = b[111:96];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5032_ = b[127:112];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5032_ = b[143:128];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5032_ = b[159:144];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5032_ = b[175:160];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5032_ = b[191:176];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5032_ = b[207:192];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5032_ = b[223:208];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5032_ = b[239:224];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5032_ = b[255:240];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5032_ = b[271:256];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5032_ = b[287:272];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5032_ = b[303:288];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5032_ = b[319:304];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5032_ = b[335:320];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5032_ = b[351:336];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5032_ = b[367:352];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5032_ = b[383:368];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5032_ = b[399:384];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5032_ = b[415:400];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5032_ = b[431:416];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5032_ = b[447:432];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5032_ = b[463:448];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5032_ = b[479:464];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5032_ = b[495:480];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5032_ = b[511:496];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5032_ = b[527:512];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5032_ = b[543:528];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5032_ = b[559:544];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5032_ = b[575:560];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5032_ = b[591:576];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5032_ = b[607:592];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5032_ = b[623:608];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5032_ = b[639:624];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5032_ = b[655:640];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5032_ = b[671:656];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5032_ = b[687:672];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5032_ = b[703:688];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5032_ = b[719:704];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5032_ = b[735:720];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5032_ = b[751:736];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5032_ = b[767:752];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5032_ = b[783:768];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5032_ = b[799:784];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5032_ = b[815:800];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5032_ = b[831:816];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5032_ = b[847:832];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5032_ = b[863:848];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5032_ = b[879:864];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5032_ = b[895:880];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5032_ = b[911:896];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5032_ = b[927:912];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5032_ = b[943:928];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5032_ = b[959:944];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5032_ = b[975:960];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5032_ = b[991:976];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5032_ = b[1007:992];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5032_ = b[1023:1008];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5032_ = b[1039:1024];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5032_ = b[1055:1040];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5032_ = b[1071:1056];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5032_ = b[1087:1072];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5032_ = b[1103:1088];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5032_ = b[1119:1104];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5032_ = b[1135:1120];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5032_ = b[1151:1136];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1167:1152];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1183:1168];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1199:1184];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1215:1200];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1231:1216];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1247:1232];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1263:1248];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1279:1264];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1295:1280];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1311:1296];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1327:1312];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1343:1328];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1359:1344];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1375:1360];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1391:1376];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1407:1392];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1423:1408];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1439:1424];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1455:1440];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1471:1456];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1487:1472];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1503:1488];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1519:1504];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1535:1520];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1551:1536];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1567:1552];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1583:1568];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1599:1584];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1615:1600];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1631:1616];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1647:1632];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1663:1648];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1679:1664];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1695:1680];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1711:1696];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1727:1712];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1743:1728];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1759:1744];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1775:1760];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1791:1776];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1807:1792];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1823:1808];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1839:1824];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1855:1840];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1871:1856];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1887:1872];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1903:1888];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1919:1904];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1935:1920];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1951:1936];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1967:1952];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1983:1968];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[1999:1984];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2015:2000];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2031:2016];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2047:2032];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2063:2048];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2079:2064];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2095:2080];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2111:2096];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2127:2112];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2143:2128];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2159:2144];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2175:2160];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2191:2176];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2207:2192];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2223:2208];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2239:2224];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2255:2240];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2271:2256];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2287:2272];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2303:2288];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2319:2304];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2335:2320];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2351:2336];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2367:2352];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2383:2368];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2399:2384];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2415:2400];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2431:2416];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2447:2432];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2463:2448];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2479:2464];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2495:2480];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2511:2496];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2527:2512];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2543:2528];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2559:2544];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2575:2560];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2591:2576];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2607:2592];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2623:2608];
      257'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2639:2624];
      257'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2655:2640];
      257'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2671:2656];
      257'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2687:2672];
      257'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2703:2688];
      257'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2719:2704];
      257'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2735:2720];
      257'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2751:2736];
      257'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2767:2752];
      257'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2783:2768];
      257'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2799:2784];
      257'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2815:2800];
      257'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2831:2816];
      257'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2847:2832];
      257'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2863:2848];
      257'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2879:2864];
      257'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2895:2880];
      257'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2911:2896];
      257'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2927:2912];
      257'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2943:2928];
      257'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2959:2944];
      257'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2975:2960];
      257'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[2991:2976];
      257'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3007:2992];
      257'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3023:3008];
      257'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3039:3024];
      257'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3055:3040];
      257'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3071:3056];
      257'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3087:3072];
      257'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3103:3088];
      257'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3119:3104];
      257'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3135:3120];
      257'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3151:3136];
      257'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3167:3152];
      257'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3183:3168];
      257'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3199:3184];
      257'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3215:3200];
      257'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3231:3216];
      257'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3247:3232];
      257'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3263:3248];
      257'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3279:3264];
      257'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3295:3280];
      257'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3311:3296];
      257'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3327:3312];
      257'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3343:3328];
      257'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3359:3344];
      257'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3375:3360];
      257'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3391:3376];
      257'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3407:3392];
      257'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3423:3408];
      257'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3439:3424];
      257'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3455:3440];
      257'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3471:3456];
      257'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3487:3472];
      257'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3503:3488];
      257'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3519:3504];
      257'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3535:3520];
      257'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3551:3536];
      257'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3567:3552];
      257'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3583:3568];
      257'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3599:3584];
      257'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3615:3600];
      257'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3631:3616];
      257'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3647:3632];
      257'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3663:3648];
      257'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3679:3664];
      257'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3695:3680];
      257'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3711:3696];
      257'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3727:3712];
      257'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3743:3728];
      257'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3759:3744];
      257'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3775:3760];
      257'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3791:3776];
      257'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3807:3792];
      257'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3823:3808];
      257'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3839:3824];
      257'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3855:3840];
      257'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3871:3856];
      257'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3887:3872];
      257'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3903:3888];
      257'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3919:3904];
      257'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3935:3920];
      257'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3951:3936];
      257'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3967:3952];
      257'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3983:3968];
      257'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[3999:3984];
      257'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4015:4000];
      257'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4031:4016];
      257'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4047:4032];
      257'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4063:4048];
      257'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4079:4064];
      257'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4095:4080];
      257'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5032_ = b[4111:4096];
      default:
        _5032_ = a;
    endcase
  endfunction
  assign lo_data0_2 = _5032_(16'b0000000000000000, { REG_lo_0, REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_, _2064_, _2063_, _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_, _1996_, _1995_, _1994_, _1993_, _1992_, _1991_, _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_ });
  assign _1938_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28367|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 9'b100000000;
  assign _1939_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28366|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111111;
  assign _1940_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28365|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111110;
  assign _1941_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28364|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111101;
  assign _1942_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28363|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111100;
  assign _1943_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28362|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111011;
  assign _1944_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28361|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111010;
  assign _1945_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28360|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111001;
  assign _1946_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28359|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11111000;
  assign _1947_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28358|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110111;
  assign _1948_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28357|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110110;
  assign _1949_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28356|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110101;
  assign _1950_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28355|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110100;
  assign _1951_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28354|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110011;
  assign _1952_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28353|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110010;
  assign _1953_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28352|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110001;
  assign _1954_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28351|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11110000;
  assign _1955_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28350|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101111;
  assign _1956_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28349|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101110;
  assign _1957_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28348|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101101;
  assign _1958_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28347|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101100;
  assign _1959_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28346|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101011;
  assign _1960_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28345|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101010;
  assign _1961_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28344|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101001;
  assign _1962_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28343|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11101000;
  assign _1963_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28342|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100111;
  assign _1964_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28341|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100110;
  assign _1965_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28340|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100101;
  assign _1966_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28339|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100100;
  assign _1967_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28338|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100011;
  assign _1968_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28337|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100010;
  assign _1969_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28336|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100001;
  assign _1970_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28335|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11100000;
  assign _1971_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28334|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011111;
  assign _1972_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28333|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011110;
  assign _1973_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28332|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011101;
  assign _1974_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28331|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011100;
  assign _1975_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28330|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011011;
  assign _1976_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28329|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011010;
  assign _1977_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28328|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011001;
  assign _1978_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28327|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11011000;
  assign _1979_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28326|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010111;
  assign _1980_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28325|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010110;
  assign _1981_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28324|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010101;
  assign _1982_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28323|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010100;
  assign _1983_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28322|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010011;
  assign _1984_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28321|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010010;
  assign _1985_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28320|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010001;
  assign _1986_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28319|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11010000;
  assign _1987_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28318|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001111;
  assign _1988_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28317|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001110;
  assign _1989_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28316|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001101;
  assign _1990_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28315|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001100;
  assign _1991_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28314|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001011;
  assign _1992_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28313|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001010;
  assign _1993_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28312|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001001;
  assign _1994_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28311|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11001000;
  assign _1995_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28310|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000111;
  assign _1996_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28309|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000110;
  assign _1997_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28308|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000101;
  assign _1998_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28307|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000100;
  assign _1999_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28306|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000011;
  assign _2000_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28305|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000010;
  assign _2001_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28304|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000001;
  assign _2002_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28303|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b11000000;
  assign _2003_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28302|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111111;
  assign _2004_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28301|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111110;
  assign _2005_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28300|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111101;
  assign _2006_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28299|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111100;
  assign _2007_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28298|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111011;
  assign _2008_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28297|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111010;
  assign _2009_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28296|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111001;
  assign _2010_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28295|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10111000;
  assign _2011_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28294|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110111;
  assign _2012_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28293|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110110;
  assign _2013_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28292|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110101;
  assign _2014_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28291|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110100;
  assign _2015_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28290|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110011;
  assign _2016_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28289|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110010;
  assign _2017_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28288|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110001;
  assign _2018_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28287|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10110000;
  assign _2019_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28286|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101111;
  assign _2020_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28285|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101110;
  assign _2021_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28284|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101101;
  assign _2022_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28283|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101100;
  assign _2023_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28282|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101011;
  assign _2024_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28281|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101010;
  assign _2025_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28280|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101001;
  assign _2026_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28279|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10101000;
  assign _2027_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28278|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100111;
  assign _2028_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28277|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100110;
  assign _2029_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28276|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100101;
  assign _2030_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28275|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100100;
  assign _2031_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28274|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100011;
  assign _2032_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28273|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100010;
  assign _2033_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28272|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100001;
  assign _2034_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28271|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10100000;
  assign _2035_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28270|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011111;
  assign _2036_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28269|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011110;
  assign _2037_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28268|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011101;
  assign _2038_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28267|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011100;
  assign _2039_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28266|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011011;
  assign _2040_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28265|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011010;
  assign _2041_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28264|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011001;
  assign _2042_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28263|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10011000;
  assign _2043_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28262|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010111;
  assign _2044_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28261|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010110;
  assign _2045_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28260|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010101;
  assign _2046_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28259|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010100;
  assign _2047_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28258|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010011;
  assign _2048_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28257|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010010;
  assign _2049_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28256|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010001;
  assign _2050_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28255|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10010000;
  assign _2051_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28254|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001111;
  assign _2052_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28253|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001110;
  assign _2053_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28252|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001101;
  assign _2054_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28251|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001100;
  assign _2055_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28250|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001011;
  assign _2056_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28249|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001010;
  assign _2057_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28248|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001001;
  assign _2058_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28247|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10001000;
  assign _2059_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28246|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000111;
  assign _2060_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28245|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000110;
  assign _2061_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28244|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000101;
  assign _2062_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28243|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000100;
  assign _2063_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28242|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000011;
  assign _2064_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28241|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000010;
  assign _2065_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28240|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000001;
  assign _2066_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28239|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 8'b10000000;
  assign _2067_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28238|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111111;
  assign _2068_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28237|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111110;
  assign _2069_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28236|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111101;
  assign _2070_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28235|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111100;
  assign _2071_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28234|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111011;
  assign _2072_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28233|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111010;
  assign _2073_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28232|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111001;
  assign _2074_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28231|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1111000;
  assign _2075_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28230|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110111;
  assign _2076_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28229|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110110;
  assign _2077_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28228|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110101;
  assign _2078_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28227|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110100;
  assign _2079_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28226|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110011;
  assign _2080_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28225|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110010;
  assign _2081_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28224|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110001;
  assign _2082_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28223|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1110000;
  assign _2083_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28222|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101111;
  assign _2084_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28221|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101110;
  assign _2085_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28220|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101101;
  assign _2086_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28219|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101100;
  assign _2087_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28218|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101011;
  assign _2088_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28217|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101010;
  assign _2089_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28216|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101001;
  assign _2090_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28215|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1101000;
  assign _2091_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28214|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100111;
  assign _2092_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28213|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100110;
  assign _2093_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28212|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100101;
  assign _2094_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28211|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100100;
  assign _2095_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28210|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100011;
  assign _2096_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28209|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100010;
  assign _2097_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28208|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100001;
  assign _2098_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28207|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1100000;
  assign _2099_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28206|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011111;
  assign _2100_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28205|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011110;
  assign _2101_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28204|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011101;
  assign _2102_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28203|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011100;
  assign _2103_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28202|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011011;
  assign _2104_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28201|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011010;
  assign _2105_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28200|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011001;
  assign _2106_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28199|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1011000;
  assign _2107_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28198|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010111;
  assign _2108_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28197|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010110;
  assign _2109_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28196|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010101;
  assign _2110_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28195|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010100;
  assign _2111_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28194|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010011;
  assign _2112_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28193|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010010;
  assign _2113_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28192|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010001;
  assign _2114_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28191|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1010000;
  assign _2115_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28190|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001111;
  assign _2116_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28189|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001110;
  assign _2117_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28188|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001101;
  assign _2118_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28187|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001100;
  assign _2119_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28186|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001011;
  assign _2120_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28185|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001010;
  assign _2121_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28184|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001001;
  assign _2122_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28183|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1001000;
  assign _2123_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28182|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000111;
  assign _2124_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28181|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000110;
  assign _2125_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28180|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000101;
  assign _2126_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28179|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000100;
  assign _2127_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28178|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000011;
  assign _2128_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28177|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000010;
  assign _2129_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28176|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000001;
  assign _2130_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28175|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 7'b1000000;
  assign _2131_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28174|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111111;
  assign _2132_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28173|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111110;
  assign _2133_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28172|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111101;
  assign _2134_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28171|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111100;
  assign _2135_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28170|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111011;
  assign _2136_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28169|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111010;
  assign _2137_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28168|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111001;
  assign _2138_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28167|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b111000;
  assign _2139_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28166|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110111;
  assign _2140_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28165|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110110;
  assign _2141_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28164|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110101;
  assign _2142_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28163|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110100;
  assign _2143_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28162|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110011;
  assign _2144_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28161|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110010;
  assign _2145_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28160|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110001;
  assign _2146_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28159|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b110000;
  assign _2147_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28158|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101111;
  assign _2148_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28157|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101110;
  assign _2149_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28156|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101101;
  assign _2150_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28155|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101100;
  assign _2151_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28154|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101011;
  assign _2152_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101010;
  assign _2153_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28152|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101001;
  assign _2154_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28151|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b101000;
  assign _2155_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28150|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100111;
  assign _2156_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28149|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100110;
  assign _2157_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28148|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100101;
  assign _2158_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28147|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100100;
  assign _2159_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28146|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100011;
  assign _2160_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28145|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100010;
  assign _2161_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28144|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100001;
  assign _2162_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28143|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 6'b100000;
  assign _2163_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28142|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11111;
  assign _2164_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28141|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11110;
  assign _2165_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28140|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11101;
  assign _2166_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28139|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11100;
  assign _2167_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28138|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11011;
  assign _2168_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28137|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11010;
  assign _2169_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11001;
  assign _2170_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28135|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b11000;
  assign _2171_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28134|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10111;
  assign _2172_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28133|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10110;
  assign _2173_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28132|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10101;
  assign _2174_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28131|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10100;
  assign _2175_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28130|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10011;
  assign _2176_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28129|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10010;
  assign _2177_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28128|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10001;
  assign _2178_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28127|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 5'b10000;
  assign _2179_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28126|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1111;
  assign _2180_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28125|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1110;
  assign _2181_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28124|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1101;
  assign _2182_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28123|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1100;
  assign _2183_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28122|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1011;
  assign _2184_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28121|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1010;
  assign _2185_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28120|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1001;
  assign _2186_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 4'b1000;
  assign _2187_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28118|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 3'b111;
  assign _2188_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28117|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 3'b110;
  assign _2189_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28116|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 3'b101;
  assign _2190_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28115|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 3'b100;
  assign _2191_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28114|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 2'b11;
  assign _2192_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28113|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 2'b10;
  assign _2193_ = p1_pipe_data[306:298] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28112|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) 1'b1;
  assign _2194_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28111|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:28110" *) p1_pipe_data[306:298];
  function [15:0] _5290_;
    input [15:0] a;
    input [4111:0] b;
    input [256:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27842|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *)
    (* parallel_case *)
    casez (s)
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5290_ = b[15:0];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5290_ = b[31:16];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5290_ = b[47:32];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5290_ = b[63:48];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5290_ = b[79:64];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5290_ = b[95:80];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5290_ = b[111:96];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5290_ = b[127:112];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5290_ = b[143:128];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5290_ = b[159:144];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5290_ = b[175:160];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5290_ = b[191:176];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5290_ = b[207:192];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5290_ = b[223:208];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5290_ = b[239:224];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5290_ = b[255:240];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5290_ = b[271:256];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5290_ = b[287:272];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5290_ = b[303:288];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5290_ = b[319:304];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5290_ = b[335:320];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5290_ = b[351:336];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5290_ = b[367:352];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5290_ = b[383:368];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5290_ = b[399:384];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5290_ = b[415:400];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5290_ = b[431:416];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5290_ = b[447:432];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5290_ = b[463:448];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5290_ = b[479:464];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5290_ = b[495:480];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5290_ = b[511:496];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5290_ = b[527:512];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5290_ = b[543:528];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5290_ = b[559:544];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5290_ = b[575:560];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5290_ = b[591:576];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5290_ = b[607:592];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5290_ = b[623:608];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5290_ = b[639:624];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5290_ = b[655:640];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5290_ = b[671:656];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5290_ = b[687:672];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5290_ = b[703:688];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5290_ = b[719:704];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5290_ = b[735:720];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5290_ = b[751:736];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5290_ = b[767:752];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5290_ = b[783:768];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5290_ = b[799:784];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5290_ = b[815:800];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5290_ = b[831:816];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5290_ = b[847:832];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5290_ = b[863:848];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5290_ = b[879:864];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5290_ = b[895:880];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5290_ = b[911:896];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5290_ = b[927:912];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5290_ = b[943:928];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5290_ = b[959:944];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5290_ = b[975:960];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5290_ = b[991:976];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5290_ = b[1007:992];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5290_ = b[1023:1008];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5290_ = b[1039:1024];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5290_ = b[1055:1040];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5290_ = b[1071:1056];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5290_ = b[1087:1072];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5290_ = b[1103:1088];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5290_ = b[1119:1104];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5290_ = b[1135:1120];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5290_ = b[1151:1136];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1167:1152];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1183:1168];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1199:1184];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1215:1200];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1231:1216];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1247:1232];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1263:1248];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1279:1264];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1295:1280];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1311:1296];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1327:1312];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1343:1328];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1359:1344];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1375:1360];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1391:1376];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1407:1392];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1423:1408];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1439:1424];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1455:1440];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1471:1456];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1487:1472];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1503:1488];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1519:1504];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1535:1520];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1551:1536];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1567:1552];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1583:1568];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1599:1584];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1615:1600];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1631:1616];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1647:1632];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1663:1648];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1679:1664];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1695:1680];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1711:1696];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1727:1712];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1743:1728];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1759:1744];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1775:1760];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1791:1776];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1807:1792];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1823:1808];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1839:1824];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1855:1840];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1871:1856];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1887:1872];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1903:1888];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1919:1904];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1935:1920];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1951:1936];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1967:1952];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1983:1968];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[1999:1984];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2015:2000];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2031:2016];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2047:2032];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2063:2048];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2079:2064];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2095:2080];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2111:2096];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2127:2112];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2143:2128];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2159:2144];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2175:2160];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2191:2176];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2207:2192];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2223:2208];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2239:2224];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2255:2240];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2271:2256];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2287:2272];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2303:2288];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2319:2304];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2335:2320];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2351:2336];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2367:2352];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2383:2368];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2399:2384];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2415:2400];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2431:2416];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2447:2432];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2463:2448];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2479:2464];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2495:2480];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2511:2496];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2527:2512];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2543:2528];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2559:2544];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2575:2560];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2591:2576];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2607:2592];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2623:2608];
      257'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2639:2624];
      257'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2655:2640];
      257'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2671:2656];
      257'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2687:2672];
      257'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2703:2688];
      257'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2719:2704];
      257'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2735:2720];
      257'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2751:2736];
      257'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2767:2752];
      257'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2783:2768];
      257'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2799:2784];
      257'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2815:2800];
      257'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2831:2816];
      257'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2847:2832];
      257'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2863:2848];
      257'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2879:2864];
      257'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2895:2880];
      257'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2911:2896];
      257'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2927:2912];
      257'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2943:2928];
      257'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2959:2944];
      257'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2975:2960];
      257'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[2991:2976];
      257'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3007:2992];
      257'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3023:3008];
      257'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3039:3024];
      257'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3055:3040];
      257'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3071:3056];
      257'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3087:3072];
      257'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3103:3088];
      257'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3119:3104];
      257'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3135:3120];
      257'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3151:3136];
      257'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3167:3152];
      257'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3183:3168];
      257'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3199:3184];
      257'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3215:3200];
      257'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3231:3216];
      257'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3247:3232];
      257'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3263:3248];
      257'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3279:3264];
      257'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3295:3280];
      257'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3311:3296];
      257'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3327:3312];
      257'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3343:3328];
      257'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3359:3344];
      257'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3375:3360];
      257'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3391:3376];
      257'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3407:3392];
      257'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3423:3408];
      257'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3439:3424];
      257'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3455:3440];
      257'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3471:3456];
      257'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3487:3472];
      257'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3503:3488];
      257'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3519:3504];
      257'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3535:3520];
      257'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3551:3536];
      257'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3567:3552];
      257'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3583:3568];
      257'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3599:3584];
      257'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3615:3600];
      257'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3631:3616];
      257'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3647:3632];
      257'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3663:3648];
      257'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3679:3664];
      257'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3695:3680];
      257'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3711:3696];
      257'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3727:3712];
      257'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3743:3728];
      257'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3759:3744];
      257'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3775:3760];
      257'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3791:3776];
      257'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3807:3792];
      257'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3823:3808];
      257'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3839:3824];
      257'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3855:3840];
      257'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3871:3856];
      257'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3887:3872];
      257'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3903:3888];
      257'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3919:3904];
      257'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3935:3920];
      257'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3951:3936];
      257'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3967:3952];
      257'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3983:3968];
      257'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[3999:3984];
      257'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4015:4000];
      257'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4031:4016];
      257'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4047:4032];
      257'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4063:4048];
      257'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4079:4064];
      257'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4095:4080];
      257'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5290_ = b[4111:4096];
      default:
        _5290_ = a;
    endcase
  endfunction
  assign lo_data0_1 = _5290_(16'b0000000000000000, { REG_lo_0, REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_, _2322_, _2321_, _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_, _2259_, _2258_, _2257_, _2256_, _2255_, _2254_, _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_ });
  assign _2195_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27842|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 9'b100000000;
  assign _2196_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27841|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111111;
  assign _2197_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27840|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111110;
  assign _2198_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27839|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111101;
  assign _2199_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27838|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111100;
  assign _2200_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27837|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111011;
  assign _2201_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27836|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111010;
  assign _2202_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27835|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111001;
  assign _2203_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27834|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11111000;
  assign _2204_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27833|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110111;
  assign _2205_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27832|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110110;
  assign _2206_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27831|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110101;
  assign _2207_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27830|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110100;
  assign _2208_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27829|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110011;
  assign _2209_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27828|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110010;
  assign _2210_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27827|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110001;
  assign _2211_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27826|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11110000;
  assign _2212_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27825|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101111;
  assign _2213_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27824|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101110;
  assign _2214_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27823|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101101;
  assign _2215_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27822|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101100;
  assign _2216_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27821|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101011;
  assign _2217_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27820|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101010;
  assign _2218_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27819|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101001;
  assign _2219_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27818|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11101000;
  assign _2220_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27817|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100111;
  assign _2221_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27816|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100110;
  assign _2222_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27815|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100101;
  assign _2223_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27814|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100100;
  assign _2224_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27813|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100011;
  assign _2225_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27812|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100010;
  assign _2226_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27811|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100001;
  assign _2227_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27810|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11100000;
  assign _2228_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27809|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011111;
  assign _2229_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27808|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011110;
  assign _2230_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27807|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011101;
  assign _2231_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27806|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011100;
  assign _2232_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27805|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011011;
  assign _2233_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27804|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011010;
  assign _2234_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27803|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011001;
  assign _2235_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27802|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11011000;
  assign _2236_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27801|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010111;
  assign _2237_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27800|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010110;
  assign _2238_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27799|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010101;
  assign _2239_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27798|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010100;
  assign _2240_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27797|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010011;
  assign _2241_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27796|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010010;
  assign _2242_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27795|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010001;
  assign _2243_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27794|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11010000;
  assign _2244_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27793|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001111;
  assign _2245_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27792|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001110;
  assign _2246_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27791|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001101;
  assign _2247_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27790|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001100;
  assign _2248_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27789|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001011;
  assign _2249_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27788|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001010;
  assign _2250_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27787|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001001;
  assign _2251_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27786|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11001000;
  assign _2252_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27785|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000111;
  assign _2253_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27784|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000110;
  assign _2254_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27783|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000101;
  assign _2255_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27782|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000100;
  assign _2256_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27781|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000011;
  assign _2257_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27780|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000010;
  assign _2258_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27779|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000001;
  assign _2259_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27778|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b11000000;
  assign _2260_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27777|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111111;
  assign _2261_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27776|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111110;
  assign _2262_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27775|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111101;
  assign _2263_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27774|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111100;
  assign _2264_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27773|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111011;
  assign _2265_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27772|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111010;
  assign _2266_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27771|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111001;
  assign _2267_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27770|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10111000;
  assign _2268_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27769|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110111;
  assign _2269_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27768|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110110;
  assign _2270_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27767|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110101;
  assign _2271_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27766|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110100;
  assign _2272_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27765|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110011;
  assign _2273_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27764|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110010;
  assign _2274_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27763|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110001;
  assign _2275_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27762|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10110000;
  assign _2276_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27761|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101111;
  assign _2277_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27760|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101110;
  assign _2278_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27759|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101101;
  assign _2279_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27758|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101100;
  assign _2280_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27757|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101011;
  assign _2281_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27756|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101010;
  assign _2282_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27755|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101001;
  assign _2283_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27754|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10101000;
  assign _2284_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27753|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100111;
  assign _2285_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27752|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100110;
  assign _2286_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27751|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100101;
  assign _2287_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27750|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100100;
  assign _2288_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27749|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100011;
  assign _2289_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27748|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100010;
  assign _2290_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27747|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100001;
  assign _2291_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27746|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10100000;
  assign _2292_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27745|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011111;
  assign _2293_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27744|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011110;
  assign _2294_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27743|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011101;
  assign _2295_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27742|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011100;
  assign _2296_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27741|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011011;
  assign _2297_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27740|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011010;
  assign _2298_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27739|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011001;
  assign _2299_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27738|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10011000;
  assign _2300_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27737|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010111;
  assign _2301_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27736|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010110;
  assign _2302_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27735|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010101;
  assign _2303_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27734|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010100;
  assign _2304_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27733|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010011;
  assign _2305_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27732|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010010;
  assign _2306_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27731|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010001;
  assign _2307_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27730|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10010000;
  assign _2308_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27729|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001111;
  assign _2309_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27728|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001110;
  assign _2310_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27727|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001101;
  assign _2311_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27726|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001100;
  assign _2312_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27725|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001011;
  assign _2313_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27724|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001010;
  assign _2314_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27723|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001001;
  assign _2315_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27722|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10001000;
  assign _2316_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27721|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000111;
  assign _2317_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27720|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000110;
  assign _2318_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27719|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000101;
  assign _2319_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27718|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000100;
  assign _2320_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27717|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000011;
  assign _2321_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27716|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000010;
  assign _2322_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27715|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000001;
  assign _2323_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27714|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 8'b10000000;
  assign _2324_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27713|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111111;
  assign _2325_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27712|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111110;
  assign _2326_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27711|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111101;
  assign _2327_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27710|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111100;
  assign _2328_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27709|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111011;
  assign _2329_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27708|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111010;
  assign _2330_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27707|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111001;
  assign _2331_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27706|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1111000;
  assign _2332_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27705|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110111;
  assign _2333_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27704|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110110;
  assign _2334_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27703|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110101;
  assign _2335_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27702|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110100;
  assign _2336_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27701|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110011;
  assign _2337_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27700|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110010;
  assign _2338_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27699|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110001;
  assign _2339_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27698|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1110000;
  assign _2340_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27697|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101111;
  assign _2341_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27696|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101110;
  assign _2342_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27695|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101101;
  assign _2343_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27694|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101100;
  assign _2344_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27693|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101011;
  assign _2345_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27692|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101010;
  assign _2346_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27691|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101001;
  assign _2347_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27690|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1101000;
  assign _2348_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27689|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100111;
  assign _2349_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27688|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100110;
  assign _2350_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27687|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100101;
  assign _2351_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27686|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100100;
  assign _2352_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27685|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100011;
  assign _2353_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27684|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100010;
  assign _2354_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27683|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100001;
  assign _2355_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27682|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1100000;
  assign _2356_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27681|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011111;
  assign _2357_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27680|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011110;
  assign _2358_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27679|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011101;
  assign _2359_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27678|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011100;
  assign _2360_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27677|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011011;
  assign _2361_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27676|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011010;
  assign _2362_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27675|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011001;
  assign _2363_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27674|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1011000;
  assign _2364_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27673|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010111;
  assign _2365_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27672|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010110;
  assign _2366_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27671|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010101;
  assign _2367_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27670|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010100;
  assign _2368_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27669|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010011;
  assign _2369_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27668|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010010;
  assign _2370_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27667|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010001;
  assign _2371_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27666|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1010000;
  assign _2372_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27665|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001111;
  assign _2373_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27664|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001110;
  assign _2374_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27663|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001101;
  assign _2375_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27662|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001100;
  assign _2376_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27661|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001011;
  assign _2377_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27660|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001010;
  assign _2378_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001001;
  assign _2379_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27658|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1001000;
  assign _2380_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27657|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000111;
  assign _2381_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27656|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000110;
  assign _2382_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27655|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000101;
  assign _2383_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27654|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000100;
  assign _2384_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27653|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000011;
  assign _2385_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27652|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000010;
  assign _2386_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27651|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000001;
  assign _2387_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27650|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 7'b1000000;
  assign _2388_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27649|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111111;
  assign _2389_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27648|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111110;
  assign _2390_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27647|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111101;
  assign _2391_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27646|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111100;
  assign _2392_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27645|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111011;
  assign _2393_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27644|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111010;
  assign _2394_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27643|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111001;
  assign _2395_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b111000;
  assign _2396_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27641|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110111;
  assign _2397_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27640|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110110;
  assign _2398_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27639|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110101;
  assign _2399_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27638|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110100;
  assign _2400_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27637|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110011;
  assign _2401_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27636|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110010;
  assign _2402_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27635|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110001;
  assign _2403_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27634|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b110000;
  assign _2404_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27633|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101111;
  assign _2405_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27632|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101110;
  assign _2406_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27631|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101101;
  assign _2407_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27630|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101100;
  assign _2408_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101011;
  assign _2409_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27628|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101010;
  assign _2410_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27627|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101001;
  assign _2411_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27626|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b101000;
  assign _2412_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27625|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100111;
  assign _2413_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27624|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100110;
  assign _2414_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27623|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100101;
  assign _2415_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27622|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100100;
  assign _2416_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27621|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100011;
  assign _2417_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27620|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100010;
  assign _2418_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27619|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100001;
  assign _2419_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27618|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 6'b100000;
  assign _2420_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27617|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11111;
  assign _2421_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27616|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11110;
  assign _2422_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27615|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11101;
  assign _2423_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27614|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11100;
  assign _2424_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27613|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11011;
  assign _2425_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11010;
  assign _2426_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27611|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11001;
  assign _2427_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27610|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b11000;
  assign _2428_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27609|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10111;
  assign _2429_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27608|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10110;
  assign _2430_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27607|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10101;
  assign _2431_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27606|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10100;
  assign _2432_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27605|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10011;
  assign _2433_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27604|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10010;
  assign _2434_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27603|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10001;
  assign _2435_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27602|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 5'b10000;
  assign _2436_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27601|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1111;
  assign _2437_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1110;
  assign _2438_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27599|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1101;
  assign _2439_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27598|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1100;
  assign _2440_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27597|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1011;
  assign _2441_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27596|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1010;
  assign _2442_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1001;
  assign _2443_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27594|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 4'b1000;
  assign _2444_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27593|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 3'b111;
  assign _2445_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27592|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 3'b110;
  assign _2446_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27591|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 3'b101;
  assign _2447_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27590|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 3'b100;
  assign _2448_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27589|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 2'b11;
  assign _2449_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27588|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 2'b10;
  assign _2450_ = p1_pipe_data[297:289] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27587|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) 1'b1;
  assign _2451_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27586|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27585" *) p1_pipe_data[297:289];
  function [15:0] _5548_;
    input [15:0] a;
    input [4111:0] b;
    input [256:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27317|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *)
    (* parallel_case *)
    casez (s)
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5548_ = b[15:0];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5548_ = b[31:16];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5548_ = b[47:32];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5548_ = b[63:48];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5548_ = b[79:64];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5548_ = b[95:80];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5548_ = b[111:96];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5548_ = b[127:112];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5548_ = b[143:128];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5548_ = b[159:144];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5548_ = b[175:160];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5548_ = b[191:176];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5548_ = b[207:192];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5548_ = b[223:208];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5548_ = b[239:224];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5548_ = b[255:240];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5548_ = b[271:256];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5548_ = b[287:272];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5548_ = b[303:288];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5548_ = b[319:304];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5548_ = b[335:320];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5548_ = b[351:336];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5548_ = b[367:352];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5548_ = b[383:368];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5548_ = b[399:384];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5548_ = b[415:400];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5548_ = b[431:416];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5548_ = b[447:432];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5548_ = b[463:448];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5548_ = b[479:464];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5548_ = b[495:480];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5548_ = b[511:496];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5548_ = b[527:512];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5548_ = b[543:528];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5548_ = b[559:544];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5548_ = b[575:560];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5548_ = b[591:576];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5548_ = b[607:592];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5548_ = b[623:608];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5548_ = b[639:624];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5548_ = b[655:640];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5548_ = b[671:656];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5548_ = b[687:672];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5548_ = b[703:688];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5548_ = b[719:704];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5548_ = b[735:720];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5548_ = b[751:736];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5548_ = b[767:752];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5548_ = b[783:768];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5548_ = b[799:784];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5548_ = b[815:800];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5548_ = b[831:816];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5548_ = b[847:832];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5548_ = b[863:848];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5548_ = b[879:864];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5548_ = b[895:880];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5548_ = b[911:896];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5548_ = b[927:912];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5548_ = b[943:928];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5548_ = b[959:944];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5548_ = b[975:960];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5548_ = b[991:976];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5548_ = b[1007:992];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5548_ = b[1023:1008];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5548_ = b[1039:1024];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5548_ = b[1055:1040];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5548_ = b[1071:1056];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5548_ = b[1087:1072];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5548_ = b[1103:1088];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5548_ = b[1119:1104];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5548_ = b[1135:1120];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5548_ = b[1151:1136];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1167:1152];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1183:1168];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1199:1184];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1215:1200];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1231:1216];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1247:1232];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1263:1248];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1279:1264];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1295:1280];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1311:1296];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1327:1312];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1343:1328];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1359:1344];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1375:1360];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1391:1376];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1407:1392];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1423:1408];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1439:1424];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1455:1440];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1471:1456];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1487:1472];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1503:1488];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1519:1504];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1535:1520];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1551:1536];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1567:1552];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1583:1568];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1599:1584];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1615:1600];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1631:1616];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1647:1632];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1663:1648];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1679:1664];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1695:1680];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1711:1696];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1727:1712];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1743:1728];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1759:1744];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1775:1760];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1791:1776];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1807:1792];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1823:1808];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1839:1824];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1855:1840];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1871:1856];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1887:1872];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1903:1888];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1919:1904];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1935:1920];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1951:1936];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1967:1952];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1983:1968];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[1999:1984];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2015:2000];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2031:2016];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2047:2032];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2063:2048];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2079:2064];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2095:2080];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2111:2096];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2127:2112];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2143:2128];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2159:2144];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2175:2160];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2191:2176];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2207:2192];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2223:2208];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2239:2224];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2255:2240];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2271:2256];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2287:2272];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2303:2288];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2319:2304];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2335:2320];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2351:2336];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2367:2352];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2383:2368];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2399:2384];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2415:2400];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2431:2416];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2447:2432];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2463:2448];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2479:2464];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2495:2480];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2511:2496];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2527:2512];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2543:2528];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2559:2544];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2575:2560];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2591:2576];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2607:2592];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2623:2608];
      257'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2639:2624];
      257'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2655:2640];
      257'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2671:2656];
      257'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2687:2672];
      257'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2703:2688];
      257'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2719:2704];
      257'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2735:2720];
      257'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2751:2736];
      257'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2767:2752];
      257'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2783:2768];
      257'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2799:2784];
      257'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2815:2800];
      257'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2831:2816];
      257'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2847:2832];
      257'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2863:2848];
      257'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2879:2864];
      257'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2895:2880];
      257'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2911:2896];
      257'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2927:2912];
      257'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2943:2928];
      257'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2959:2944];
      257'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2975:2960];
      257'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[2991:2976];
      257'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3007:2992];
      257'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3023:3008];
      257'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3039:3024];
      257'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3055:3040];
      257'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3071:3056];
      257'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3087:3072];
      257'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3103:3088];
      257'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3119:3104];
      257'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3135:3120];
      257'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3151:3136];
      257'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3167:3152];
      257'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3183:3168];
      257'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3199:3184];
      257'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3215:3200];
      257'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3231:3216];
      257'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3247:3232];
      257'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3263:3248];
      257'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3279:3264];
      257'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3295:3280];
      257'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3311:3296];
      257'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3327:3312];
      257'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3343:3328];
      257'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3359:3344];
      257'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3375:3360];
      257'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3391:3376];
      257'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3407:3392];
      257'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3423:3408];
      257'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3439:3424];
      257'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3455:3440];
      257'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3471:3456];
      257'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3487:3472];
      257'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3503:3488];
      257'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3519:3504];
      257'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3535:3520];
      257'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3551:3536];
      257'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3567:3552];
      257'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3583:3568];
      257'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3599:3584];
      257'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3615:3600];
      257'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3631:3616];
      257'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3647:3632];
      257'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3663:3648];
      257'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3679:3664];
      257'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3695:3680];
      257'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3711:3696];
      257'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3727:3712];
      257'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3743:3728];
      257'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3759:3744];
      257'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3775:3760];
      257'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3791:3776];
      257'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3807:3792];
      257'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3823:3808];
      257'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3839:3824];
      257'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3855:3840];
      257'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3871:3856];
      257'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3887:3872];
      257'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3903:3888];
      257'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3919:3904];
      257'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3935:3920];
      257'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3951:3936];
      257'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3967:3952];
      257'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3983:3968];
      257'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[3999:3984];
      257'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4015:4000];
      257'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4031:4016];
      257'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4047:4032];
      257'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4063:4048];
      257'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4079:4064];
      257'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4095:4080];
      257'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5548_ = b[4111:4096];
      default:
        _5548_ = a;
    endcase
  endfunction
  assign lo_data0_0 = _5548_(16'b0000000000000000, { REG_lo_0, REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_, _2580_, _2579_, _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_, _2522_, _2521_, _2520_, _2519_, _2518_, _2517_, _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_ });
  assign _2452_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27317|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 9'b100000000;
  assign _2453_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27316|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111111;
  assign _2454_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27315|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111110;
  assign _2455_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27314|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111101;
  assign _2456_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27313|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111100;
  assign _2457_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27312|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111011;
  assign _2458_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27311|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111010;
  assign _2459_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27310|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111001;
  assign _2460_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27309|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11111000;
  assign _2461_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27308|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110111;
  assign _2462_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27307|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110110;
  assign _2463_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27306|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110101;
  assign _2464_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27305|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110100;
  assign _2465_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27304|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110011;
  assign _2466_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27303|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110010;
  assign _2467_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27302|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110001;
  assign _2468_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27301|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11110000;
  assign _2469_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27300|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101111;
  assign _2470_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27299|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101110;
  assign _2471_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27298|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101101;
  assign _2472_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27297|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101100;
  assign _2473_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27296|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101011;
  assign _2474_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27295|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101010;
  assign _2475_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27294|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101001;
  assign _2476_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27293|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11101000;
  assign _2477_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27292|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100111;
  assign _2478_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27291|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100110;
  assign _2479_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27290|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100101;
  assign _2480_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27289|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100100;
  assign _2481_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27288|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100011;
  assign _2482_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27287|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100010;
  assign _2483_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27286|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100001;
  assign _2484_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27285|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11100000;
  assign _2485_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27284|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011111;
  assign _2486_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27283|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011110;
  assign _2487_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27282|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011101;
  assign _2488_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27281|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011100;
  assign _2489_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27280|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011011;
  assign _2490_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27279|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011010;
  assign _2491_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27278|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011001;
  assign _2492_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27277|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11011000;
  assign _2493_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27276|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010111;
  assign _2494_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27275|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010110;
  assign _2495_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27274|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010101;
  assign _2496_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27273|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010100;
  assign _2497_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27272|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010011;
  assign _2498_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27271|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010010;
  assign _2499_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27270|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010001;
  assign _2500_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27269|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11010000;
  assign _2501_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27268|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001111;
  assign _2502_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27267|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001110;
  assign _2503_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27266|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001101;
  assign _2504_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27265|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001100;
  assign _2505_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27264|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001011;
  assign _2506_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27263|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001010;
  assign _2507_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27262|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001001;
  assign _2508_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27261|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11001000;
  assign _2509_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27260|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000111;
  assign _2510_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27259|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000110;
  assign _2511_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27258|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000101;
  assign _2512_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27257|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000100;
  assign _2513_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27256|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000011;
  assign _2514_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27255|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000010;
  assign _2515_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27254|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000001;
  assign _2516_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27253|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b11000000;
  assign _2517_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27252|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111111;
  assign _2518_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27251|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111110;
  assign _2519_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27250|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111101;
  assign _2520_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27249|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111100;
  assign _2521_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27248|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111011;
  assign _2522_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27247|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111010;
  assign _2523_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27246|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111001;
  assign _2524_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27245|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10111000;
  assign _2525_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27244|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110111;
  assign _2526_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27243|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110110;
  assign _2527_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27242|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110101;
  assign _2528_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27241|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110100;
  assign _2529_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27240|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110011;
  assign _2530_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27239|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110010;
  assign _2531_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27238|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110001;
  assign _2532_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27237|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10110000;
  assign _2533_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27236|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101111;
  assign _2534_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27235|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101110;
  assign _2535_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27234|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101101;
  assign _2536_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27233|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101100;
  assign _2537_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27232|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101011;
  assign _2538_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27231|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101010;
  assign _2539_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27230|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101001;
  assign _2540_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27229|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10101000;
  assign _2541_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27228|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100111;
  assign _2542_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27227|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100110;
  assign _2543_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27226|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100101;
  assign _2544_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27225|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100100;
  assign _2545_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27224|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100011;
  assign _2546_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27223|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100010;
  assign _2547_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27222|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100001;
  assign _2548_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27221|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10100000;
  assign _2549_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27220|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011111;
  assign _2550_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27219|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011110;
  assign _2551_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27218|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011101;
  assign _2552_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27217|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011100;
  assign _2553_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27216|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011011;
  assign _2554_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27215|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011010;
  assign _2555_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27214|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011001;
  assign _2556_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27213|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10011000;
  assign _2557_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27212|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010111;
  assign _2558_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27211|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010110;
  assign _2559_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27210|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010101;
  assign _2560_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27209|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010100;
  assign _2561_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27208|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010011;
  assign _2562_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27207|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010010;
  assign _2563_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27206|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010001;
  assign _2564_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27205|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10010000;
  assign _2565_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27204|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001111;
  assign _2566_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27203|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001110;
  assign _2567_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27202|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001101;
  assign _2568_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27201|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001100;
  assign _2569_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27200|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001011;
  assign _2570_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27199|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001010;
  assign _2571_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27198|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001001;
  assign _2572_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27197|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10001000;
  assign _2573_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27196|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000111;
  assign _2574_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27195|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000110;
  assign _2575_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27194|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000101;
  assign _2576_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27193|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000100;
  assign _2577_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27192|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000011;
  assign _2578_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27191|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000010;
  assign _2579_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27190|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000001;
  assign _2580_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27189|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 8'b10000000;
  assign _2581_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27188|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111111;
  assign _2582_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27187|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111110;
  assign _2583_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27186|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111101;
  assign _2584_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27185|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111100;
  assign _2585_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27184|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111011;
  assign _2586_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27183|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111010;
  assign _2587_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27182|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111001;
  assign _2588_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27181|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1111000;
  assign _2589_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27180|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110111;
  assign _2590_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27179|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110110;
  assign _2591_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27178|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110101;
  assign _2592_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27177|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110100;
  assign _2593_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27176|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110011;
  assign _2594_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27175|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110010;
  assign _2595_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27174|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110001;
  assign _2596_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27173|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1110000;
  assign _2597_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27172|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101111;
  assign _2598_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27171|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101110;
  assign _2599_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27170|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101101;
  assign _2600_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27169|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101100;
  assign _2601_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27168|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101011;
  assign _2602_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27167|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101010;
  assign _2603_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27166|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101001;
  assign _2604_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27165|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1101000;
  assign _2605_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27164|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100111;
  assign _2606_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27163|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100110;
  assign _2607_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27162|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100101;
  assign _2608_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27161|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100100;
  assign _2609_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27160|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100011;
  assign _2610_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27159|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100010;
  assign _2611_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27158|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100001;
  assign _2612_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27157|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1100000;
  assign _2613_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27156|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011111;
  assign _2614_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27155|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011110;
  assign _2615_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27154|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011101;
  assign _2616_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011100;
  assign _2617_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27152|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011011;
  assign _2618_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27151|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011010;
  assign _2619_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27150|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011001;
  assign _2620_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27149|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1011000;
  assign _2621_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27148|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010111;
  assign _2622_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27147|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010110;
  assign _2623_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27146|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010101;
  assign _2624_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27145|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010100;
  assign _2625_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27144|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010011;
  assign _2626_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27143|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010010;
  assign _2627_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27142|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010001;
  assign _2628_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27141|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1010000;
  assign _2629_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27140|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001111;
  assign _2630_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27139|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001110;
  assign _2631_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27138|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001101;
  assign _2632_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27137|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001100;
  assign _2633_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001011;
  assign _2634_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27135|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001010;
  assign _2635_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27134|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001001;
  assign _2636_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27133|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1001000;
  assign _2637_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27132|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000111;
  assign _2638_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27131|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000110;
  assign _2639_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27130|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000101;
  assign _2640_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27129|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000100;
  assign _2641_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27128|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000011;
  assign _2642_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27127|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000010;
  assign _2643_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27126|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000001;
  assign _2644_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27125|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 7'b1000000;
  assign _2645_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27124|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111111;
  assign _2646_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27123|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111110;
  assign _2647_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27122|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111101;
  assign _2648_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27121|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111100;
  assign _2649_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27120|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111011;
  assign _2650_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111010;
  assign _2651_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27118|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111001;
  assign _2652_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27117|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b111000;
  assign _2653_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27116|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110111;
  assign _2654_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27115|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110110;
  assign _2655_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27114|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110101;
  assign _2656_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27113|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110100;
  assign _2657_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27112|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110011;
  assign _2658_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27111|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110010;
  assign _2659_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27110|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110001;
  assign _2660_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27109|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b110000;
  assign _2661_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27108|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101111;
  assign _2662_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27107|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101110;
  assign _2663_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27106|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101101;
  assign _2664_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27105|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101100;
  assign _2665_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27104|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101011;
  assign _2666_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27103|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101010;
  assign _2667_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27102|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101001;
  assign _2668_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27101|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b101000;
  assign _2669_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27100|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100111;
  assign _2670_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27099|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100110;
  assign _2671_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27098|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100101;
  assign _2672_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27097|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100100;
  assign _2673_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27096|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100011;
  assign _2674_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27095|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100010;
  assign _2675_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27094|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100001;
  assign _2676_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27093|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 6'b100000;
  assign _2677_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27092|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11111;
  assign _2678_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27091|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11110;
  assign _2679_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27090|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11101;
  assign _2680_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27089|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11100;
  assign _2681_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27088|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11011;
  assign _2682_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27087|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11010;
  assign _2683_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27086|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11001;
  assign _2684_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27085|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b11000;
  assign _2685_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27084|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10111;
  assign _2686_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27083|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10110;
  assign _2687_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27082|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10101;
  assign _2688_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27081|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10100;
  assign _2689_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27080|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10011;
  assign _2690_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27079|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10010;
  assign _2691_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27078|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10001;
  assign _2692_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27077|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 5'b10000;
  assign _2693_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27076|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1111;
  assign _2694_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27075|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1110;
  assign _2695_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27074|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1101;
  assign _2696_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27073|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1100;
  assign _2697_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27072|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1011;
  assign _2698_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27071|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1010;
  assign _2699_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27070|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1001;
  assign _2700_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27069|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 4'b1000;
  assign _2701_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27068|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 3'b111;
  assign _2702_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27067|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 3'b110;
  assign _2703_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27066|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 3'b101;
  assign _2704_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27065|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 3'b100;
  assign _2705_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27064|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 2'b11;
  assign _2706_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27063|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 2'b10;
  assign _2707_ = p1_pipe_data[288:280] == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27062|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) 1'b1;
  assign _2708_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27061|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:27060" *) p1_pipe_data[288:280];
  function [15:0] _5806_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:26792|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:26536" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _5806_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _5806_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _5806_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _5806_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _5806_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _5806_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _5806_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _5806_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _5806_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _5806_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _5806_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _5806_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _5806_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _5806_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _5806_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _5806_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _5806_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _5806_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _5806_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _5806_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _5806_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _5806_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _5806_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _5806_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _5806_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _5806_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _5806_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _5806_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _5806_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _5806_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _5806_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _5806_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _5806_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _5806_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _5806_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _5806_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _5806_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _5806_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _5806_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _5806_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _5806_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _5806_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _5806_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _5806_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _5806_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _5806_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _5806_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _5806_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _5806_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _5806_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _5806_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _5806_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _5806_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _5806_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _5806_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _5806_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _5806_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _5806_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _5806_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _5806_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _5806_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _5806_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _5806_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _5806_ = b[1023:1008];
      default:
        _5806_ = a;
    endcase
  endfunction
  assign le_data1_3 = _5806_(16'b0000000000000000, { REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_ });
  function [15:0] _5807_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:26269|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:26013" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _5807_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _5807_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _5807_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _5807_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _5807_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _5807_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _5807_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _5807_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _5807_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _5807_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _5807_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _5807_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _5807_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _5807_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _5807_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _5807_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _5807_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _5807_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _5807_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _5807_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _5807_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _5807_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _5807_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _5807_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _5807_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _5807_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _5807_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _5807_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _5807_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _5807_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _5807_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _5807_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _5807_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _5807_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _5807_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _5807_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _5807_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _5807_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _5807_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _5807_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _5807_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _5807_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _5807_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _5807_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _5807_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _5807_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _5807_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _5807_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _5807_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _5807_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _5807_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _5807_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _5807_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _5807_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _5807_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _5807_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _5807_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _5807_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _5807_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _5807_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _5807_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _5807_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _5807_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _5807_ = b[1023:1008];
      default:
        _5807_ = a;
    endcase
  endfunction
  assign le_data1_2 = _5807_(16'b0000000000000000, { REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_ });
  function [15:0] _5808_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:25746|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:25490" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _5808_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _5808_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _5808_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _5808_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _5808_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _5808_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _5808_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _5808_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _5808_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _5808_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _5808_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _5808_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _5808_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _5808_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _5808_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _5808_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _5808_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _5808_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _5808_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _5808_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _5808_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _5808_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _5808_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _5808_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _5808_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _5808_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _5808_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _5808_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _5808_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _5808_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _5808_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _5808_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _5808_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _5808_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _5808_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _5808_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _5808_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _5808_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _5808_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _5808_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _5808_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _5808_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _5808_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _5808_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _5808_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _5808_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _5808_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _5808_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _5808_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _5808_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _5808_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _5808_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _5808_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _5808_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _5808_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _5808_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _5808_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _5808_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _5808_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _5808_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _5808_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _5808_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _5808_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _5808_ = b[1023:1008];
      default:
        _5808_ = a;
    endcase
  endfunction
  assign le_data1_1 = _5808_(16'b0000000000000000, { REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_ });
  function [15:0] _5809_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:25223|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:24967" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _5809_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _5809_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _5809_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _5809_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _5809_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _5809_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _5809_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _5809_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _5809_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _5809_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _5809_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _5809_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _5809_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _5809_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _5809_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _5809_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _5809_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _5809_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _5809_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _5809_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _5809_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _5809_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _5809_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _5809_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _5809_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _5809_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _5809_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _5809_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _5809_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _5809_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _5809_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _5809_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _5809_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _5809_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _5809_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _5809_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _5809_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _5809_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _5809_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _5809_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _5809_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _5809_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _5809_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _5809_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _5809_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _5809_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _5809_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _5809_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _5809_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _5809_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _5809_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _5809_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _5809_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _5809_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _5809_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _5809_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _5809_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _5809_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _5809_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _5809_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _5809_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _5809_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _5809_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _5809_ = b[1023:1008];
      default:
        _5809_ = a;
    endcase
  endfunction
  assign le_data1_0 = _5809_(16'b0000000000000000, { REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_ });
  function [15:0] _5810_;
    input [15:0] a;
    input [1039:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:24700|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:24443" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _5810_ = b[15:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _5810_ = b[31:16];
      65'b??????????????????????????????????????????????????????????????1??:
        _5810_ = b[47:32];
      65'b?????????????????????????????????????????????????????????????1???:
        _5810_ = b[63:48];
      65'b????????????????????????????????????????????????????????????1????:
        _5810_ = b[79:64];
      65'b???????????????????????????????????????????????????????????1?????:
        _5810_ = b[95:80];
      65'b??????????????????????????????????????????????????????????1??????:
        _5810_ = b[111:96];
      65'b?????????????????????????????????????????????????????????1???????:
        _5810_ = b[127:112];
      65'b????????????????????????????????????????????????????????1????????:
        _5810_ = b[143:128];
      65'b???????????????????????????????????????????????????????1?????????:
        _5810_ = b[159:144];
      65'b??????????????????????????????????????????????????????1??????????:
        _5810_ = b[175:160];
      65'b?????????????????????????????????????????????????????1???????????:
        _5810_ = b[191:176];
      65'b????????????????????????????????????????????????????1????????????:
        _5810_ = b[207:192];
      65'b???????????????????????????????????????????????????1?????????????:
        _5810_ = b[223:208];
      65'b??????????????????????????????????????????????????1??????????????:
        _5810_ = b[239:224];
      65'b?????????????????????????????????????????????????1???????????????:
        _5810_ = b[255:240];
      65'b????????????????????????????????????????????????1????????????????:
        _5810_ = b[271:256];
      65'b???????????????????????????????????????????????1?????????????????:
        _5810_ = b[287:272];
      65'b??????????????????????????????????????????????1??????????????????:
        _5810_ = b[303:288];
      65'b?????????????????????????????????????????????1???????????????????:
        _5810_ = b[319:304];
      65'b????????????????????????????????????????????1????????????????????:
        _5810_ = b[335:320];
      65'b???????????????????????????????????????????1?????????????????????:
        _5810_ = b[351:336];
      65'b??????????????????????????????????????????1??????????????????????:
        _5810_ = b[367:352];
      65'b?????????????????????????????????????????1???????????????????????:
        _5810_ = b[383:368];
      65'b????????????????????????????????????????1????????????????????????:
        _5810_ = b[399:384];
      65'b???????????????????????????????????????1?????????????????????????:
        _5810_ = b[415:400];
      65'b??????????????????????????????????????1??????????????????????????:
        _5810_ = b[431:416];
      65'b?????????????????????????????????????1???????????????????????????:
        _5810_ = b[447:432];
      65'b????????????????????????????????????1????????????????????????????:
        _5810_ = b[463:448];
      65'b???????????????????????????????????1?????????????????????????????:
        _5810_ = b[479:464];
      65'b??????????????????????????????????1??????????????????????????????:
        _5810_ = b[495:480];
      65'b?????????????????????????????????1???????????????????????????????:
        _5810_ = b[511:496];
      65'b????????????????????????????????1????????????????????????????????:
        _5810_ = b[527:512];
      65'b???????????????????????????????1?????????????????????????????????:
        _5810_ = b[543:528];
      65'b??????????????????????????????1??????????????????????????????????:
        _5810_ = b[559:544];
      65'b?????????????????????????????1???????????????????????????????????:
        _5810_ = b[575:560];
      65'b????????????????????????????1????????????????????????????????????:
        _5810_ = b[591:576];
      65'b???????????????????????????1?????????????????????????????????????:
        _5810_ = b[607:592];
      65'b??????????????????????????1??????????????????????????????????????:
        _5810_ = b[623:608];
      65'b?????????????????????????1???????????????????????????????????????:
        _5810_ = b[639:624];
      65'b????????????????????????1????????????????????????????????????????:
        _5810_ = b[655:640];
      65'b???????????????????????1?????????????????????????????????????????:
        _5810_ = b[671:656];
      65'b??????????????????????1??????????????????????????????????????????:
        _5810_ = b[687:672];
      65'b?????????????????????1???????????????????????????????????????????:
        _5810_ = b[703:688];
      65'b????????????????????1????????????????????????????????????????????:
        _5810_ = b[719:704];
      65'b???????????????????1?????????????????????????????????????????????:
        _5810_ = b[735:720];
      65'b??????????????????1??????????????????????????????????????????????:
        _5810_ = b[751:736];
      65'b?????????????????1???????????????????????????????????????????????:
        _5810_ = b[767:752];
      65'b????????????????1????????????????????????????????????????????????:
        _5810_ = b[783:768];
      65'b???????????????1?????????????????????????????????????????????????:
        _5810_ = b[799:784];
      65'b??????????????1??????????????????????????????????????????????????:
        _5810_ = b[815:800];
      65'b?????????????1???????????????????????????????????????????????????:
        _5810_ = b[831:816];
      65'b????????????1????????????????????????????????????????????????????:
        _5810_ = b[847:832];
      65'b???????????1?????????????????????????????????????????????????????:
        _5810_ = b[863:848];
      65'b??????????1??????????????????????????????????????????????????????:
        _5810_ = b[879:864];
      65'b?????????1???????????????????????????????????????????????????????:
        _5810_ = b[895:880];
      65'b????????1????????????????????????????????????????????????????????:
        _5810_ = b[911:896];
      65'b???????1?????????????????????????????????????????????????????????:
        _5810_ = b[927:912];
      65'b??????1??????????????????????????????????????????????????????????:
        _5810_ = b[943:928];
      65'b?????1???????????????????????????????????????????????????????????:
        _5810_ = b[959:944];
      65'b????1????????????????????????????????????????????????????????????:
        _5810_ = b[975:960];
      65'b???1?????????????????????????????????????????????????????????????:
        _5810_ = b[991:976];
      65'b??1??????????????????????????????????????????????????????????????:
        _5810_ = b[1007:992];
      65'b?1???????????????????????????????????????????????????????????????:
        _5810_ = b[1023:1008];
      65'b1????????????????????????????????????????????????????????????????:
        _5810_ = b[1039:1024];
      default:
        _5810_ = a;
    endcase
  endfunction
  assign le_data0_3 = _5810_(16'b0000000000000000, { REG_le_0, REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_ });
  function [15:0] _5811_;
    input [15:0] a;
    input [1039:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:24175|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:23918" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _5811_ = b[15:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _5811_ = b[31:16];
      65'b??????????????????????????????????????????????????????????????1??:
        _5811_ = b[47:32];
      65'b?????????????????????????????????????????????????????????????1???:
        _5811_ = b[63:48];
      65'b????????????????????????????????????????????????????????????1????:
        _5811_ = b[79:64];
      65'b???????????????????????????????????????????????????????????1?????:
        _5811_ = b[95:80];
      65'b??????????????????????????????????????????????????????????1??????:
        _5811_ = b[111:96];
      65'b?????????????????????????????????????????????????????????1???????:
        _5811_ = b[127:112];
      65'b????????????????????????????????????????????????????????1????????:
        _5811_ = b[143:128];
      65'b???????????????????????????????????????????????????????1?????????:
        _5811_ = b[159:144];
      65'b??????????????????????????????????????????????????????1??????????:
        _5811_ = b[175:160];
      65'b?????????????????????????????????????????????????????1???????????:
        _5811_ = b[191:176];
      65'b????????????????????????????????????????????????????1????????????:
        _5811_ = b[207:192];
      65'b???????????????????????????????????????????????????1?????????????:
        _5811_ = b[223:208];
      65'b??????????????????????????????????????????????????1??????????????:
        _5811_ = b[239:224];
      65'b?????????????????????????????????????????????????1???????????????:
        _5811_ = b[255:240];
      65'b????????????????????????????????????????????????1????????????????:
        _5811_ = b[271:256];
      65'b???????????????????????????????????????????????1?????????????????:
        _5811_ = b[287:272];
      65'b??????????????????????????????????????????????1??????????????????:
        _5811_ = b[303:288];
      65'b?????????????????????????????????????????????1???????????????????:
        _5811_ = b[319:304];
      65'b????????????????????????????????????????????1????????????????????:
        _5811_ = b[335:320];
      65'b???????????????????????????????????????????1?????????????????????:
        _5811_ = b[351:336];
      65'b??????????????????????????????????????????1??????????????????????:
        _5811_ = b[367:352];
      65'b?????????????????????????????????????????1???????????????????????:
        _5811_ = b[383:368];
      65'b????????????????????????????????????????1????????????????????????:
        _5811_ = b[399:384];
      65'b???????????????????????????????????????1?????????????????????????:
        _5811_ = b[415:400];
      65'b??????????????????????????????????????1??????????????????????????:
        _5811_ = b[431:416];
      65'b?????????????????????????????????????1???????????????????????????:
        _5811_ = b[447:432];
      65'b????????????????????????????????????1????????????????????????????:
        _5811_ = b[463:448];
      65'b???????????????????????????????????1?????????????????????????????:
        _5811_ = b[479:464];
      65'b??????????????????????????????????1??????????????????????????????:
        _5811_ = b[495:480];
      65'b?????????????????????????????????1???????????????????????????????:
        _5811_ = b[511:496];
      65'b????????????????????????????????1????????????????????????????????:
        _5811_ = b[527:512];
      65'b???????????????????????????????1?????????????????????????????????:
        _5811_ = b[543:528];
      65'b??????????????????????????????1??????????????????????????????????:
        _5811_ = b[559:544];
      65'b?????????????????????????????1???????????????????????????????????:
        _5811_ = b[575:560];
      65'b????????????????????????????1????????????????????????????????????:
        _5811_ = b[591:576];
      65'b???????????????????????????1?????????????????????????????????????:
        _5811_ = b[607:592];
      65'b??????????????????????????1??????????????????????????????????????:
        _5811_ = b[623:608];
      65'b?????????????????????????1???????????????????????????????????????:
        _5811_ = b[639:624];
      65'b????????????????????????1????????????????????????????????????????:
        _5811_ = b[655:640];
      65'b???????????????????????1?????????????????????????????????????????:
        _5811_ = b[671:656];
      65'b??????????????????????1??????????????????????????????????????????:
        _5811_ = b[687:672];
      65'b?????????????????????1???????????????????????????????????????????:
        _5811_ = b[703:688];
      65'b????????????????????1????????????????????????????????????????????:
        _5811_ = b[719:704];
      65'b???????????????????1?????????????????????????????????????????????:
        _5811_ = b[735:720];
      65'b??????????????????1??????????????????????????????????????????????:
        _5811_ = b[751:736];
      65'b?????????????????1???????????????????????????????????????????????:
        _5811_ = b[767:752];
      65'b????????????????1????????????????????????????????????????????????:
        _5811_ = b[783:768];
      65'b???????????????1?????????????????????????????????????????????????:
        _5811_ = b[799:784];
      65'b??????????????1??????????????????????????????????????????????????:
        _5811_ = b[815:800];
      65'b?????????????1???????????????????????????????????????????????????:
        _5811_ = b[831:816];
      65'b????????????1????????????????????????????????????????????????????:
        _5811_ = b[847:832];
      65'b???????????1?????????????????????????????????????????????????????:
        _5811_ = b[863:848];
      65'b??????????1??????????????????????????????????????????????????????:
        _5811_ = b[879:864];
      65'b?????????1???????????????????????????????????????????????????????:
        _5811_ = b[895:880];
      65'b????????1????????????????????????????????????????????????????????:
        _5811_ = b[911:896];
      65'b???????1?????????????????????????????????????????????????????????:
        _5811_ = b[927:912];
      65'b??????1??????????????????????????????????????????????????????????:
        _5811_ = b[943:928];
      65'b?????1???????????????????????????????????????????????????????????:
        _5811_ = b[959:944];
      65'b????1????????????????????????????????????????????????????????????:
        _5811_ = b[975:960];
      65'b???1?????????????????????????????????????????????????????????????:
        _5811_ = b[991:976];
      65'b??1??????????????????????????????????????????????????????????????:
        _5811_ = b[1007:992];
      65'b?1???????????????????????????????????????????????????????????????:
        _5811_ = b[1023:1008];
      65'b1????????????????????????????????????????????????????????????????:
        _5811_ = b[1039:1024];
      default:
        _5811_ = a;
    endcase
  endfunction
  assign le_data0_2 = _5811_(16'b0000000000000000, { REG_le_0, REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_ });
  function [15:0] _5812_;
    input [15:0] a;
    input [1039:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:23650|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:23393" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _5812_ = b[15:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _5812_ = b[31:16];
      65'b??????????????????????????????????????????????????????????????1??:
        _5812_ = b[47:32];
      65'b?????????????????????????????????????????????????????????????1???:
        _5812_ = b[63:48];
      65'b????????????????????????????????????????????????????????????1????:
        _5812_ = b[79:64];
      65'b???????????????????????????????????????????????????????????1?????:
        _5812_ = b[95:80];
      65'b??????????????????????????????????????????????????????????1??????:
        _5812_ = b[111:96];
      65'b?????????????????????????????????????????????????????????1???????:
        _5812_ = b[127:112];
      65'b????????????????????????????????????????????????????????1????????:
        _5812_ = b[143:128];
      65'b???????????????????????????????????????????????????????1?????????:
        _5812_ = b[159:144];
      65'b??????????????????????????????????????????????????????1??????????:
        _5812_ = b[175:160];
      65'b?????????????????????????????????????????????????????1???????????:
        _5812_ = b[191:176];
      65'b????????????????????????????????????????????????????1????????????:
        _5812_ = b[207:192];
      65'b???????????????????????????????????????????????????1?????????????:
        _5812_ = b[223:208];
      65'b??????????????????????????????????????????????????1??????????????:
        _5812_ = b[239:224];
      65'b?????????????????????????????????????????????????1???????????????:
        _5812_ = b[255:240];
      65'b????????????????????????????????????????????????1????????????????:
        _5812_ = b[271:256];
      65'b???????????????????????????????????????????????1?????????????????:
        _5812_ = b[287:272];
      65'b??????????????????????????????????????????????1??????????????????:
        _5812_ = b[303:288];
      65'b?????????????????????????????????????????????1???????????????????:
        _5812_ = b[319:304];
      65'b????????????????????????????????????????????1????????????????????:
        _5812_ = b[335:320];
      65'b???????????????????????????????????????????1?????????????????????:
        _5812_ = b[351:336];
      65'b??????????????????????????????????????????1??????????????????????:
        _5812_ = b[367:352];
      65'b?????????????????????????????????????????1???????????????????????:
        _5812_ = b[383:368];
      65'b????????????????????????????????????????1????????????????????????:
        _5812_ = b[399:384];
      65'b???????????????????????????????????????1?????????????????????????:
        _5812_ = b[415:400];
      65'b??????????????????????????????????????1??????????????????????????:
        _5812_ = b[431:416];
      65'b?????????????????????????????????????1???????????????????????????:
        _5812_ = b[447:432];
      65'b????????????????????????????????????1????????????????????????????:
        _5812_ = b[463:448];
      65'b???????????????????????????????????1?????????????????????????????:
        _5812_ = b[479:464];
      65'b??????????????????????????????????1??????????????????????????????:
        _5812_ = b[495:480];
      65'b?????????????????????????????????1???????????????????????????????:
        _5812_ = b[511:496];
      65'b????????????????????????????????1????????????????????????????????:
        _5812_ = b[527:512];
      65'b???????????????????????????????1?????????????????????????????????:
        _5812_ = b[543:528];
      65'b??????????????????????????????1??????????????????????????????????:
        _5812_ = b[559:544];
      65'b?????????????????????????????1???????????????????????????????????:
        _5812_ = b[575:560];
      65'b????????????????????????????1????????????????????????????????????:
        _5812_ = b[591:576];
      65'b???????????????????????????1?????????????????????????????????????:
        _5812_ = b[607:592];
      65'b??????????????????????????1??????????????????????????????????????:
        _5812_ = b[623:608];
      65'b?????????????????????????1???????????????????????????????????????:
        _5812_ = b[639:624];
      65'b????????????????????????1????????????????????????????????????????:
        _5812_ = b[655:640];
      65'b???????????????????????1?????????????????????????????????????????:
        _5812_ = b[671:656];
      65'b??????????????????????1??????????????????????????????????????????:
        _5812_ = b[687:672];
      65'b?????????????????????1???????????????????????????????????????????:
        _5812_ = b[703:688];
      65'b????????????????????1????????????????????????????????????????????:
        _5812_ = b[719:704];
      65'b???????????????????1?????????????????????????????????????????????:
        _5812_ = b[735:720];
      65'b??????????????????1??????????????????????????????????????????????:
        _5812_ = b[751:736];
      65'b?????????????????1???????????????????????????????????????????????:
        _5812_ = b[767:752];
      65'b????????????????1????????????????????????????????????????????????:
        _5812_ = b[783:768];
      65'b???????????????1?????????????????????????????????????????????????:
        _5812_ = b[799:784];
      65'b??????????????1??????????????????????????????????????????????????:
        _5812_ = b[815:800];
      65'b?????????????1???????????????????????????????????????????????????:
        _5812_ = b[831:816];
      65'b????????????1????????????????????????????????????????????????????:
        _5812_ = b[847:832];
      65'b???????????1?????????????????????????????????????????????????????:
        _5812_ = b[863:848];
      65'b??????????1??????????????????????????????????????????????????????:
        _5812_ = b[879:864];
      65'b?????????1???????????????????????????????????????????????????????:
        _5812_ = b[895:880];
      65'b????????1????????????????????????????????????????????????????????:
        _5812_ = b[911:896];
      65'b???????1?????????????????????????????????????????????????????????:
        _5812_ = b[927:912];
      65'b??????1??????????????????????????????????????????????????????????:
        _5812_ = b[943:928];
      65'b?????1???????????????????????????????????????????????????????????:
        _5812_ = b[959:944];
      65'b????1????????????????????????????????????????????????????????????:
        _5812_ = b[975:960];
      65'b???1?????????????????????????????????????????????????????????????:
        _5812_ = b[991:976];
      65'b??1??????????????????????????????????????????????????????????????:
        _5812_ = b[1007:992];
      65'b?1???????????????????????????????????????????????????????????????:
        _5812_ = b[1023:1008];
      65'b1????????????????????????????????????????????????????????????????:
        _5812_ = b[1039:1024];
      default:
        _5812_ = a;
    endcase
  endfunction
  assign le_data0_1 = _5812_(16'b0000000000000000, { REG_le_0, REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_ });
  function [15:0] _5813_;
    input [15:0] a;
    input [1039:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:23125|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22868" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _5813_ = b[15:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _5813_ = b[31:16];
      65'b??????????????????????????????????????????????????????????????1??:
        _5813_ = b[47:32];
      65'b?????????????????????????????????????????????????????????????1???:
        _5813_ = b[63:48];
      65'b????????????????????????????????????????????????????????????1????:
        _5813_ = b[79:64];
      65'b???????????????????????????????????????????????????????????1?????:
        _5813_ = b[95:80];
      65'b??????????????????????????????????????????????????????????1??????:
        _5813_ = b[111:96];
      65'b?????????????????????????????????????????????????????????1???????:
        _5813_ = b[127:112];
      65'b????????????????????????????????????????????????????????1????????:
        _5813_ = b[143:128];
      65'b???????????????????????????????????????????????????????1?????????:
        _5813_ = b[159:144];
      65'b??????????????????????????????????????????????????????1??????????:
        _5813_ = b[175:160];
      65'b?????????????????????????????????????????????????????1???????????:
        _5813_ = b[191:176];
      65'b????????????????????????????????????????????????????1????????????:
        _5813_ = b[207:192];
      65'b???????????????????????????????????????????????????1?????????????:
        _5813_ = b[223:208];
      65'b??????????????????????????????????????????????????1??????????????:
        _5813_ = b[239:224];
      65'b?????????????????????????????????????????????????1???????????????:
        _5813_ = b[255:240];
      65'b????????????????????????????????????????????????1????????????????:
        _5813_ = b[271:256];
      65'b???????????????????????????????????????????????1?????????????????:
        _5813_ = b[287:272];
      65'b??????????????????????????????????????????????1??????????????????:
        _5813_ = b[303:288];
      65'b?????????????????????????????????????????????1???????????????????:
        _5813_ = b[319:304];
      65'b????????????????????????????????????????????1????????????????????:
        _5813_ = b[335:320];
      65'b???????????????????????????????????????????1?????????????????????:
        _5813_ = b[351:336];
      65'b??????????????????????????????????????????1??????????????????????:
        _5813_ = b[367:352];
      65'b?????????????????????????????????????????1???????????????????????:
        _5813_ = b[383:368];
      65'b????????????????????????????????????????1????????????????????????:
        _5813_ = b[399:384];
      65'b???????????????????????????????????????1?????????????????????????:
        _5813_ = b[415:400];
      65'b??????????????????????????????????????1??????????????????????????:
        _5813_ = b[431:416];
      65'b?????????????????????????????????????1???????????????????????????:
        _5813_ = b[447:432];
      65'b????????????????????????????????????1????????????????????????????:
        _5813_ = b[463:448];
      65'b???????????????????????????????????1?????????????????????????????:
        _5813_ = b[479:464];
      65'b??????????????????????????????????1??????????????????????????????:
        _5813_ = b[495:480];
      65'b?????????????????????????????????1???????????????????????????????:
        _5813_ = b[511:496];
      65'b????????????????????????????????1????????????????????????????????:
        _5813_ = b[527:512];
      65'b???????????????????????????????1?????????????????????????????????:
        _5813_ = b[543:528];
      65'b??????????????????????????????1??????????????????????????????????:
        _5813_ = b[559:544];
      65'b?????????????????????????????1???????????????????????????????????:
        _5813_ = b[575:560];
      65'b????????????????????????????1????????????????????????????????????:
        _5813_ = b[591:576];
      65'b???????????????????????????1?????????????????????????????????????:
        _5813_ = b[607:592];
      65'b??????????????????????????1??????????????????????????????????????:
        _5813_ = b[623:608];
      65'b?????????????????????????1???????????????????????????????????????:
        _5813_ = b[639:624];
      65'b????????????????????????1????????????????????????????????????????:
        _5813_ = b[655:640];
      65'b???????????????????????1?????????????????????????????????????????:
        _5813_ = b[671:656];
      65'b??????????????????????1??????????????????????????????????????????:
        _5813_ = b[687:672];
      65'b?????????????????????1???????????????????????????????????????????:
        _5813_ = b[703:688];
      65'b????????????????????1????????????????????????????????????????????:
        _5813_ = b[719:704];
      65'b???????????????????1?????????????????????????????????????????????:
        _5813_ = b[735:720];
      65'b??????????????????1??????????????????????????????????????????????:
        _5813_ = b[751:736];
      65'b?????????????????1???????????????????????????????????????????????:
        _5813_ = b[767:752];
      65'b????????????????1????????????????????????????????????????????????:
        _5813_ = b[783:768];
      65'b???????????????1?????????????????????????????????????????????????:
        _5813_ = b[799:784];
      65'b??????????????1??????????????????????????????????????????????????:
        _5813_ = b[815:800];
      65'b?????????????1???????????????????????????????????????????????????:
        _5813_ = b[831:816];
      65'b????????????1????????????????????????????????????????????????????:
        _5813_ = b[847:832];
      65'b???????????1?????????????????????????????????????????????????????:
        _5813_ = b[863:848];
      65'b??????????1??????????????????????????????????????????????????????:
        _5813_ = b[879:864];
      65'b?????????1???????????????????????????????????????????????????????:
        _5813_ = b[895:880];
      65'b????????1????????????????????????????????????????????????????????:
        _5813_ = b[911:896];
      65'b???????1?????????????????????????????????????????????????????????:
        _5813_ = b[927:912];
      65'b??????1??????????????????????????????????????????????????????????:
        _5813_ = b[943:928];
      65'b?????1???????????????????????????????????????????????????????????:
        _5813_ = b[959:944];
      65'b????1????????????????????????????????????????????????????????????:
        _5813_ = b[975:960];
      65'b???1?????????????????????????????????????????????????????????????:
        _5813_ = b[991:976];
      65'b??1??????????????????????????????????????????????????????????????:
        _5813_ = b[1007:992];
      65'b?1???????????????????????????????????????????????????????????????:
        _5813_ = b[1023:1008];
      65'b1????????????????????????????????????????????????????????????????:
        _5813_ = b[1039:1024];
      default:
        _5813_ = a;
    endcase
  endfunction
  assign le_data0_0 = _5813_(16'b0000000000000000, { REG_le_0, REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_ });
  assign _0331_ = reg2dp_perf_lut_en ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22587" *) perf_lut_lo_hit_cnt_nxt : perf_lut_lo_hit_cnt_cur;
  assign _0330_ = reg2dp_perf_lut_en ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22544" *) perf_lut_le_hit_cnt_nxt : perf_lut_le_hit_cnt_cur;
  assign _0329_ = reg2dp_perf_lut_en ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22501" *) perf_lut_hybrid_cnt_nxt : perf_lut_hybrid_cnt_cur;
  assign _0333_ = reg2dp_perf_lut_en ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22454" *) perf_lut_uflow_cnt_nxt : perf_lut_uflow_cnt_cur;
  assign _0332_ = reg2dp_perf_lut_en ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22411" *) perf_lut_oflow_cnt_nxt : perf_lut_oflow_cnt_cur;
  assign _0238_ = lo_wr_en_256 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21965" *) reg2dp_lut_int_data : REG_lo_256;
  assign _0237_ = lo_wr_en_255 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21903" *) reg2dp_lut_int_data : REG_lo_255;
  assign _0236_ = lo_wr_en_254 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21841" *) reg2dp_lut_int_data : REG_lo_254;
  assign _0235_ = lo_wr_en_253 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21779" *) reg2dp_lut_int_data : REG_lo_253;
  assign _0234_ = lo_wr_en_252 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21717" *) reg2dp_lut_int_data : REG_lo_252;
  assign _0233_ = lo_wr_en_251 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21655" *) reg2dp_lut_int_data : REG_lo_251;
  assign _0232_ = lo_wr_en_250 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21593" *) reg2dp_lut_int_data : REG_lo_250;
  assign _0230_ = lo_wr_en_249 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21531" *) reg2dp_lut_int_data : REG_lo_249;
  assign _0229_ = lo_wr_en_248 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21469" *) reg2dp_lut_int_data : REG_lo_248;
  assign _0228_ = lo_wr_en_247 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21407" *) reg2dp_lut_int_data : REG_lo_247;
  assign _0227_ = lo_wr_en_246 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21345" *) reg2dp_lut_int_data : REG_lo_246;
  assign _0226_ = lo_wr_en_245 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21283" *) reg2dp_lut_int_data : REG_lo_245;
  assign _0225_ = lo_wr_en_244 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21221" *) reg2dp_lut_int_data : REG_lo_244;
  assign _0224_ = lo_wr_en_243 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21159" *) reg2dp_lut_int_data : REG_lo_243;
  assign _0223_ = lo_wr_en_242 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21097" *) reg2dp_lut_int_data : REG_lo_242;
  assign _0222_ = lo_wr_en_241 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:21035" *) reg2dp_lut_int_data : REG_lo_241;
  assign _0221_ = lo_wr_en_240 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20973" *) reg2dp_lut_int_data : REG_lo_240;
  assign _0219_ = lo_wr_en_239 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20911" *) reg2dp_lut_int_data : REG_lo_239;
  assign _0218_ = lo_wr_en_238 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20849" *) reg2dp_lut_int_data : REG_lo_238;
  assign _0217_ = lo_wr_en_237 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20787" *) reg2dp_lut_int_data : REG_lo_237;
  assign _0216_ = lo_wr_en_236 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20725" *) reg2dp_lut_int_data : REG_lo_236;
  assign _0215_ = lo_wr_en_235 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20663" *) reg2dp_lut_int_data : REG_lo_235;
  assign _0214_ = lo_wr_en_234 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20601" *) reg2dp_lut_int_data : REG_lo_234;
  assign _0213_ = lo_wr_en_233 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20539" *) reg2dp_lut_int_data : REG_lo_233;
  assign _0212_ = lo_wr_en_232 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20477" *) reg2dp_lut_int_data : REG_lo_232;
  assign _0211_ = lo_wr_en_231 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20415" *) reg2dp_lut_int_data : REG_lo_231;
  assign _0210_ = lo_wr_en_230 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20353" *) reg2dp_lut_int_data : REG_lo_230;
  assign _0208_ = lo_wr_en_229 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20291" *) reg2dp_lut_int_data : REG_lo_229;
  assign _0207_ = lo_wr_en_228 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20229" *) reg2dp_lut_int_data : REG_lo_228;
  assign _0206_ = lo_wr_en_227 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20167" *) reg2dp_lut_int_data : REG_lo_227;
  assign _0205_ = lo_wr_en_226 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20105" *) reg2dp_lut_int_data : REG_lo_226;
  assign _0204_ = lo_wr_en_225 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:20043" *) reg2dp_lut_int_data : REG_lo_225;
  assign _0203_ = lo_wr_en_224 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19981" *) reg2dp_lut_int_data : REG_lo_224;
  assign _0202_ = lo_wr_en_223 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19919" *) reg2dp_lut_int_data : REG_lo_223;
  assign _0201_ = lo_wr_en_222 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19857" *) reg2dp_lut_int_data : REG_lo_222;
  assign _0200_ = lo_wr_en_221 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19795" *) reg2dp_lut_int_data : REG_lo_221;
  assign _0199_ = lo_wr_en_220 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19733" *) reg2dp_lut_int_data : REG_lo_220;
  assign _0197_ = lo_wr_en_219 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19671" *) reg2dp_lut_int_data : REG_lo_219;
  assign _0196_ = lo_wr_en_218 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19609" *) reg2dp_lut_int_data : REG_lo_218;
  assign _0195_ = lo_wr_en_217 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19547" *) reg2dp_lut_int_data : REG_lo_217;
  assign _0194_ = lo_wr_en_216 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19485" *) reg2dp_lut_int_data : REG_lo_216;
  assign _0193_ = lo_wr_en_215 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19423" *) reg2dp_lut_int_data : REG_lo_215;
  assign _0192_ = lo_wr_en_214 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19361" *) reg2dp_lut_int_data : REG_lo_214;
  assign _0191_ = lo_wr_en_213 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19299" *) reg2dp_lut_int_data : REG_lo_213;
  assign _0190_ = lo_wr_en_212 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19237" *) reg2dp_lut_int_data : REG_lo_212;
  assign _0189_ = lo_wr_en_211 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19175" *) reg2dp_lut_int_data : REG_lo_211;
  assign _0188_ = lo_wr_en_210 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19113" *) reg2dp_lut_int_data : REG_lo_210;
  assign _0186_ = lo_wr_en_209 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:19051" *) reg2dp_lut_int_data : REG_lo_209;
  assign _0185_ = lo_wr_en_208 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18989" *) reg2dp_lut_int_data : REG_lo_208;
  assign _0184_ = lo_wr_en_207 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18927" *) reg2dp_lut_int_data : REG_lo_207;
  assign _0183_ = lo_wr_en_206 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18865" *) reg2dp_lut_int_data : REG_lo_206;
  assign _0182_ = lo_wr_en_205 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18803" *) reg2dp_lut_int_data : REG_lo_205;
  assign _0181_ = lo_wr_en_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18741" *) reg2dp_lut_int_data : REG_lo_204;
  assign _0180_ = lo_wr_en_203 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18679" *) reg2dp_lut_int_data : REG_lo_203;
  assign _0179_ = lo_wr_en_202 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18617" *) reg2dp_lut_int_data : REG_lo_202;
  assign _0178_ = lo_wr_en_201 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18555" *) reg2dp_lut_int_data : REG_lo_201;
  assign _0177_ = lo_wr_en_200 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18493" *) reg2dp_lut_int_data : REG_lo_200;
  assign _0174_ = lo_wr_en_199 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18431" *) reg2dp_lut_int_data : REG_lo_199;
  assign _0173_ = lo_wr_en_198 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18369" *) reg2dp_lut_int_data : REG_lo_198;
  assign _0172_ = lo_wr_en_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18307" *) reg2dp_lut_int_data : REG_lo_197;
  assign _0171_ = lo_wr_en_196 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18245" *) reg2dp_lut_int_data : REG_lo_196;
  assign _0170_ = lo_wr_en_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18183" *) reg2dp_lut_int_data : REG_lo_195;
  assign _0169_ = lo_wr_en_194 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18121" *) reg2dp_lut_int_data : REG_lo_194;
  assign _0168_ = lo_wr_en_193 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:18059" *) reg2dp_lut_int_data : REG_lo_193;
  assign _0167_ = lo_wr_en_192 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17997" *) reg2dp_lut_int_data : REG_lo_192;
  assign _0166_ = lo_wr_en_191 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17935" *) reg2dp_lut_int_data : REG_lo_191;
  assign _0165_ = lo_wr_en_190 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17873" *) reg2dp_lut_int_data : REG_lo_190;
  assign _0163_ = lo_wr_en_189 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17811" *) reg2dp_lut_int_data : REG_lo_189;
  assign _0162_ = lo_wr_en_188 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17749" *) reg2dp_lut_int_data : REG_lo_188;
  assign _0161_ = lo_wr_en_187 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17687" *) reg2dp_lut_int_data : REG_lo_187;
  assign _0160_ = lo_wr_en_186 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17625" *) reg2dp_lut_int_data : REG_lo_186;
  assign _0159_ = lo_wr_en_185 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17563" *) reg2dp_lut_int_data : REG_lo_185;
  assign _0158_ = lo_wr_en_184 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17501" *) reg2dp_lut_int_data : REG_lo_184;
  assign _0157_ = lo_wr_en_183 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17439" *) reg2dp_lut_int_data : REG_lo_183;
  assign _0156_ = lo_wr_en_182 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17377" *) reg2dp_lut_int_data : REG_lo_182;
  assign _0155_ = lo_wr_en_181 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17315" *) reg2dp_lut_int_data : REG_lo_181;
  assign _0154_ = lo_wr_en_180 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17253" *) reg2dp_lut_int_data : REG_lo_180;
  assign _0152_ = lo_wr_en_179 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17191" *) reg2dp_lut_int_data : REG_lo_179;
  assign _0151_ = lo_wr_en_178 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17129" *) reg2dp_lut_int_data : REG_lo_178;
  assign _0150_ = lo_wr_en_177 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17067" *) reg2dp_lut_int_data : REG_lo_177;
  assign _0149_ = lo_wr_en_176 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:17005" *) reg2dp_lut_int_data : REG_lo_176;
  assign _0148_ = lo_wr_en_175 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16943" *) reg2dp_lut_int_data : REG_lo_175;
  assign _0147_ = lo_wr_en_174 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16881" *) reg2dp_lut_int_data : REG_lo_174;
  assign _0146_ = lo_wr_en_173 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16819" *) reg2dp_lut_int_data : REG_lo_173;
  assign _0145_ = lo_wr_en_172 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16757" *) reg2dp_lut_int_data : REG_lo_172;
  assign _0144_ = lo_wr_en_171 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16695" *) reg2dp_lut_int_data : REG_lo_171;
  assign _0143_ = lo_wr_en_170 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16633" *) reg2dp_lut_int_data : REG_lo_170;
  assign _0141_ = lo_wr_en_169 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16571" *) reg2dp_lut_int_data : REG_lo_169;
  assign _0140_ = lo_wr_en_168 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16509" *) reg2dp_lut_int_data : REG_lo_168;
  assign _0139_ = lo_wr_en_167 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16447" *) reg2dp_lut_int_data : REG_lo_167;
  assign _0138_ = lo_wr_en_166 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16385" *) reg2dp_lut_int_data : REG_lo_166;
  assign _0137_ = lo_wr_en_165 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16323" *) reg2dp_lut_int_data : REG_lo_165;
  assign _0136_ = lo_wr_en_164 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16261" *) reg2dp_lut_int_data : REG_lo_164;
  assign _0135_ = lo_wr_en_163 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16199" *) reg2dp_lut_int_data : REG_lo_163;
  assign _0134_ = lo_wr_en_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16137" *) reg2dp_lut_int_data : REG_lo_162;
  assign _0133_ = lo_wr_en_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16075" *) reg2dp_lut_int_data : REG_lo_161;
  assign _0132_ = lo_wr_en_160 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:16013" *) reg2dp_lut_int_data : REG_lo_160;
  assign _0130_ = lo_wr_en_159 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15951" *) reg2dp_lut_int_data : REG_lo_159;
  assign _0129_ = lo_wr_en_158 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15889" *) reg2dp_lut_int_data : REG_lo_158;
  assign _0128_ = lo_wr_en_157 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15827" *) reg2dp_lut_int_data : REG_lo_157;
  assign _0127_ = lo_wr_en_156 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15765" *) reg2dp_lut_int_data : REG_lo_156;
  assign _0126_ = lo_wr_en_155 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15703" *) reg2dp_lut_int_data : REG_lo_155;
  assign _0125_ = lo_wr_en_154 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15641" *) reg2dp_lut_int_data : REG_lo_154;
  assign _0124_ = lo_wr_en_153 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15579" *) reg2dp_lut_int_data : REG_lo_153;
  assign _0123_ = lo_wr_en_152 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15517" *) reg2dp_lut_int_data : REG_lo_152;
  assign _0122_ = lo_wr_en_151 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15455" *) reg2dp_lut_int_data : REG_lo_151;
  assign _0121_ = lo_wr_en_150 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15393" *) reg2dp_lut_int_data : REG_lo_150;
  assign _0119_ = lo_wr_en_149 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15331" *) reg2dp_lut_int_data : REG_lo_149;
  assign _0118_ = lo_wr_en_148 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15269" *) reg2dp_lut_int_data : REG_lo_148;
  assign _0117_ = lo_wr_en_147 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15207" *) reg2dp_lut_int_data : REG_lo_147;
  assign _0116_ = lo_wr_en_146 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15145" *) reg2dp_lut_int_data : REG_lo_146;
  assign _0115_ = lo_wr_en_145 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15083" *) reg2dp_lut_int_data : REG_lo_145;
  assign _0114_ = lo_wr_en_144 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:15021" *) reg2dp_lut_int_data : REG_lo_144;
  assign _0113_ = lo_wr_en_143 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14959" *) reg2dp_lut_int_data : REG_lo_143;
  assign _0112_ = lo_wr_en_142 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14897" *) reg2dp_lut_int_data : REG_lo_142;
  assign _0111_ = lo_wr_en_141 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14835" *) reg2dp_lut_int_data : REG_lo_141;
  assign _0110_ = lo_wr_en_140 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14773" *) reg2dp_lut_int_data : REG_lo_140;
  assign _0108_ = lo_wr_en_139 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14711" *) reg2dp_lut_int_data : REG_lo_139;
  assign _0107_ = lo_wr_en_138 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14649" *) reg2dp_lut_int_data : REG_lo_138;
  assign _0106_ = lo_wr_en_137 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14587" *) reg2dp_lut_int_data : REG_lo_137;
  assign _0105_ = lo_wr_en_136 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14525" *) reg2dp_lut_int_data : REG_lo_136;
  assign _0104_ = lo_wr_en_135 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14463" *) reg2dp_lut_int_data : REG_lo_135;
  assign _0103_ = lo_wr_en_134 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14401" *) reg2dp_lut_int_data : REG_lo_134;
  assign _0102_ = lo_wr_en_133 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14339" *) reg2dp_lut_int_data : REG_lo_133;
  assign _0101_ = lo_wr_en_132 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14277" *) reg2dp_lut_int_data : REG_lo_132;
  assign _0100_ = lo_wr_en_131 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14215" *) reg2dp_lut_int_data : REG_lo_131;
  assign _0099_ = lo_wr_en_130 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14153" *) reg2dp_lut_int_data : REG_lo_130;
  assign _0097_ = lo_wr_en_129 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14091" *) reg2dp_lut_int_data : REG_lo_129;
  assign _0096_ = lo_wr_en_128 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:14029" *) reg2dp_lut_int_data : REG_lo_128;
  assign _0095_ = lo_wr_en_127 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13967" *) reg2dp_lut_int_data : REG_lo_127;
  assign _0094_ = lo_wr_en_126 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13905" *) reg2dp_lut_int_data : REG_lo_126;
  assign _0093_ = lo_wr_en_125 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13843" *) reg2dp_lut_int_data : REG_lo_125;
  assign _0092_ = lo_wr_en_124 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13781" *) reg2dp_lut_int_data : REG_lo_124;
  assign _0091_ = lo_wr_en_123 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13719" *) reg2dp_lut_int_data : REG_lo_123;
  assign _0090_ = lo_wr_en_122 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13657" *) reg2dp_lut_int_data : REG_lo_122;
  assign _0089_ = lo_wr_en_121 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13595" *) reg2dp_lut_int_data : REG_lo_121;
  assign _0088_ = lo_wr_en_120 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13533" *) reg2dp_lut_int_data : REG_lo_120;
  assign _0086_ = lo_wr_en_119 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13471" *) reg2dp_lut_int_data : REG_lo_119;
  assign _0085_ = lo_wr_en_118 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13409" *) reg2dp_lut_int_data : REG_lo_118;
  assign _0084_ = lo_wr_en_117 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13347" *) reg2dp_lut_int_data : REG_lo_117;
  assign _0083_ = lo_wr_en_116 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13285" *) reg2dp_lut_int_data : REG_lo_116;
  assign _0082_ = lo_wr_en_115 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13223" *) reg2dp_lut_int_data : REG_lo_115;
  assign _0081_ = lo_wr_en_114 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13161" *) reg2dp_lut_int_data : REG_lo_114;
  assign _0080_ = lo_wr_en_113 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13099" *) reg2dp_lut_int_data : REG_lo_113;
  assign _0079_ = lo_wr_en_112 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:13037" *) reg2dp_lut_int_data : REG_lo_112;
  assign _0078_ = lo_wr_en_111 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12975" *) reg2dp_lut_int_data : REG_lo_111;
  assign _0077_ = lo_wr_en_110 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12913" *) reg2dp_lut_int_data : REG_lo_110;
  assign _0075_ = lo_wr_en_109 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12851" *) reg2dp_lut_int_data : REG_lo_109;
  assign _0074_ = lo_wr_en_108 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12789" *) reg2dp_lut_int_data : REG_lo_108;
  assign _0073_ = lo_wr_en_107 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12727" *) reg2dp_lut_int_data : REG_lo_107;
  assign _0072_ = lo_wr_en_106 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12665" *) reg2dp_lut_int_data : REG_lo_106;
  assign _0071_ = lo_wr_en_105 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12603" *) reg2dp_lut_int_data : REG_lo_105;
  assign _0070_ = lo_wr_en_104 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12541" *) reg2dp_lut_int_data : REG_lo_104;
  assign _0069_ = lo_wr_en_103 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12479" *) reg2dp_lut_int_data : REG_lo_103;
  assign _0068_ = lo_wr_en_102 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12417" *) reg2dp_lut_int_data : REG_lo_102;
  assign _0067_ = lo_wr_en_101 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12355" *) reg2dp_lut_int_data : REG_lo_101;
  assign _0066_ = lo_wr_en_100 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12293" *) reg2dp_lut_int_data : REG_lo_100;
  assign _0320_ = lo_wr_en_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12231" *) reg2dp_lut_int_data : REG_lo_99;
  assign _0319_ = lo_wr_en_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12169" *) reg2dp_lut_int_data : REG_lo_98;
  assign _0318_ = lo_wr_en_97 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12107" *) reg2dp_lut_int_data : REG_lo_97;
  assign _0317_ = lo_wr_en_96 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:12045" *) reg2dp_lut_int_data : REG_lo_96;
  assign _0316_ = lo_wr_en_95 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11983" *) reg2dp_lut_int_data : REG_lo_95;
  assign _0315_ = lo_wr_en_94 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11921" *) reg2dp_lut_int_data : REG_lo_94;
  assign _0314_ = lo_wr_en_93 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11859" *) reg2dp_lut_int_data : REG_lo_93;
  assign _0313_ = lo_wr_en_92 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11797" *) reg2dp_lut_int_data : REG_lo_92;
  assign _0312_ = lo_wr_en_91 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11735" *) reg2dp_lut_int_data : REG_lo_91;
  assign _0311_ = lo_wr_en_90 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11673" *) reg2dp_lut_int_data : REG_lo_90;
  assign _0309_ = lo_wr_en_89 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11611" *) reg2dp_lut_int_data : REG_lo_89;
  assign _0308_ = lo_wr_en_88 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11549" *) reg2dp_lut_int_data : REG_lo_88;
  assign _0307_ = lo_wr_en_87 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11487" *) reg2dp_lut_int_data : REG_lo_87;
  assign _0306_ = lo_wr_en_86 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11425" *) reg2dp_lut_int_data : REG_lo_86;
  assign _0305_ = lo_wr_en_85 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11363" *) reg2dp_lut_int_data : REG_lo_85;
  assign _0304_ = lo_wr_en_84 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11301" *) reg2dp_lut_int_data : REG_lo_84;
  assign _0303_ = lo_wr_en_83 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11239" *) reg2dp_lut_int_data : REG_lo_83;
  assign _0302_ = lo_wr_en_82 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11177" *) reg2dp_lut_int_data : REG_lo_82;
  assign _0301_ = lo_wr_en_81 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11115" *) reg2dp_lut_int_data : REG_lo_81;
  assign _0300_ = lo_wr_en_80 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:11053" *) reg2dp_lut_int_data : REG_lo_80;
  assign _0298_ = lo_wr_en_79 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10991" *) reg2dp_lut_int_data : REG_lo_79;
  assign _0297_ = lo_wr_en_78 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10929" *) reg2dp_lut_int_data : REG_lo_78;
  assign _0296_ = lo_wr_en_77 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10867" *) reg2dp_lut_int_data : REG_lo_77;
  assign _0295_ = lo_wr_en_76 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10805" *) reg2dp_lut_int_data : REG_lo_76;
  assign _0294_ = lo_wr_en_75 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10743" *) reg2dp_lut_int_data : REG_lo_75;
  assign _0293_ = lo_wr_en_74 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10681" *) reg2dp_lut_int_data : REG_lo_74;
  assign _0292_ = lo_wr_en_73 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10619" *) reg2dp_lut_int_data : REG_lo_73;
  assign _0291_ = lo_wr_en_72 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10557" *) reg2dp_lut_int_data : REG_lo_72;
  assign _0290_ = lo_wr_en_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10495" *) reg2dp_lut_int_data : REG_lo_71;
  assign _0289_ = lo_wr_en_70 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10433" *) reg2dp_lut_int_data : REG_lo_70;
  assign _0287_ = lo_wr_en_69 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10371" *) reg2dp_lut_int_data : REG_lo_69;
  assign _0286_ = lo_wr_en_68 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10309" *) reg2dp_lut_int_data : REG_lo_68;
  assign _0285_ = lo_wr_en_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10247" *) reg2dp_lut_int_data : REG_lo_67;
  assign _0284_ = lo_wr_en_66 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10185" *) reg2dp_lut_int_data : REG_lo_66;
  assign _0283_ = lo_wr_en_65 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10123" *) reg2dp_lut_int_data : REG_lo_65;
  assign _0282_ = lo_wr_en_64 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:10061" *) reg2dp_lut_int_data : REG_lo_64;
  assign _0281_ = lo_wr_en_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9999" *) reg2dp_lut_int_data : REG_lo_63;
  assign _0280_ = lo_wr_en_62 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9937" *) reg2dp_lut_int_data : REG_lo_62;
  assign _0279_ = lo_wr_en_61 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9875" *) reg2dp_lut_int_data : REG_lo_61;
  assign _0278_ = lo_wr_en_60 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9813" *) reg2dp_lut_int_data : REG_lo_60;
  assign _0276_ = lo_wr_en_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9751" *) reg2dp_lut_int_data : REG_lo_59;
  assign _0275_ = lo_wr_en_58 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9689" *) reg2dp_lut_int_data : REG_lo_58;
  assign _0274_ = lo_wr_en_57 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9627" *) reg2dp_lut_int_data : REG_lo_57;
  assign _0273_ = lo_wr_en_56 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9565" *) reg2dp_lut_int_data : REG_lo_56;
  assign _0272_ = lo_wr_en_55 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9503" *) reg2dp_lut_int_data : REG_lo_55;
  assign _0271_ = lo_wr_en_54 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9441" *) reg2dp_lut_int_data : REG_lo_54;
  assign _0270_ = lo_wr_en_53 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9379" *) reg2dp_lut_int_data : REG_lo_53;
  assign _0269_ = lo_wr_en_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9317" *) reg2dp_lut_int_data : REG_lo_52;
  assign _0268_ = lo_wr_en_51 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9255" *) reg2dp_lut_int_data : REG_lo_51;
  assign _0267_ = lo_wr_en_50 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9193" *) reg2dp_lut_int_data : REG_lo_50;
  assign _0265_ = lo_wr_en_49 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9131" *) reg2dp_lut_int_data : REG_lo_49;
  assign _0264_ = lo_wr_en_48 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9069" *) reg2dp_lut_int_data : REG_lo_48;
  assign _0263_ = lo_wr_en_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:9007" *) reg2dp_lut_int_data : REG_lo_47;
  assign _0262_ = lo_wr_en_46 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8945" *) reg2dp_lut_int_data : REG_lo_46;
  assign _0261_ = lo_wr_en_45 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8883" *) reg2dp_lut_int_data : REG_lo_45;
  assign _0260_ = lo_wr_en_44 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8821" *) reg2dp_lut_int_data : REG_lo_44;
  assign _0259_ = lo_wr_en_43 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8759" *) reg2dp_lut_int_data : REG_lo_43;
  assign _0258_ = lo_wr_en_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8697" *) reg2dp_lut_int_data : REG_lo_42;
  assign _0257_ = lo_wr_en_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8635" *) reg2dp_lut_int_data : REG_lo_41;
  assign _0256_ = lo_wr_en_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8573" *) reg2dp_lut_int_data : REG_lo_40;
  assign _0254_ = lo_wr_en_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8511" *) reg2dp_lut_int_data : REG_lo_39;
  assign _0253_ = lo_wr_en_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8449" *) reg2dp_lut_int_data : REG_lo_38;
  assign _0252_ = lo_wr_en_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8387" *) reg2dp_lut_int_data : REG_lo_37;
  assign _0251_ = lo_wr_en_36 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8325" *) reg2dp_lut_int_data : REG_lo_36;
  assign _0250_ = lo_wr_en_35 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8263" *) reg2dp_lut_int_data : REG_lo_35;
  assign _0249_ = lo_wr_en_34 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8201" *) reg2dp_lut_int_data : REG_lo_34;
  assign _0248_ = lo_wr_en_33 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8139" *) reg2dp_lut_int_data : REG_lo_33;
  assign _0247_ = lo_wr_en_32 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8077" *) reg2dp_lut_int_data : REG_lo_32;
  assign _0246_ = lo_wr_en_31 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:8015" *) reg2dp_lut_int_data : REG_lo_31;
  assign _0245_ = lo_wr_en_30 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7953" *) reg2dp_lut_int_data : REG_lo_30;
  assign _0243_ = lo_wr_en_29 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7891" *) reg2dp_lut_int_data : REG_lo_29;
  assign _0242_ = lo_wr_en_28 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7829" *) reg2dp_lut_int_data : REG_lo_28;
  assign _0241_ = lo_wr_en_27 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7767" *) reg2dp_lut_int_data : REG_lo_27;
  assign _0240_ = lo_wr_en_26 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7705" *) reg2dp_lut_int_data : REG_lo_26;
  assign _0239_ = lo_wr_en_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7643" *) reg2dp_lut_int_data : REG_lo_25;
  assign _0231_ = lo_wr_en_24 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7581" *) reg2dp_lut_int_data : REG_lo_24;
  assign _0220_ = lo_wr_en_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7519" *) reg2dp_lut_int_data : REG_lo_23;
  assign _0209_ = lo_wr_en_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7457" *) reg2dp_lut_int_data : REG_lo_22;
  assign _0198_ = lo_wr_en_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7395" *) reg2dp_lut_int_data : REG_lo_21;
  assign _0187_ = lo_wr_en_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7333" *) reg2dp_lut_int_data : REG_lo_20;
  assign _0175_ = lo_wr_en_19 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7271" *) reg2dp_lut_int_data : REG_lo_19;
  assign _0164_ = lo_wr_en_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7209" *) reg2dp_lut_int_data : REG_lo_18;
  assign _0153_ = lo_wr_en_17 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7147" *) reg2dp_lut_int_data : REG_lo_17;
  assign _0142_ = lo_wr_en_16 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7085" *) reg2dp_lut_int_data : REG_lo_16;
  assign _0131_ = lo_wr_en_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:7023" *) reg2dp_lut_int_data : REG_lo_15;
  assign _0120_ = lo_wr_en_14 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6961" *) reg2dp_lut_int_data : REG_lo_14;
  assign _0109_ = lo_wr_en_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6899" *) reg2dp_lut_int_data : REG_lo_13;
  assign _0098_ = lo_wr_en_12 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6837" *) reg2dp_lut_int_data : REG_lo_12;
  assign _0087_ = lo_wr_en_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6775" *) reg2dp_lut_int_data : REG_lo_11;
  assign _0076_ = lo_wr_en_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6713" *) reg2dp_lut_int_data : REG_lo_10;
  assign _0321_ = lo_wr_en_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6651" *) reg2dp_lut_int_data : REG_lo_9;
  assign _0310_ = lo_wr_en_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6589" *) reg2dp_lut_int_data : REG_lo_8;
  assign _0299_ = lo_wr_en_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6527" *) reg2dp_lut_int_data : REG_lo_7;
  assign _0288_ = lo_wr_en_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6465" *) reg2dp_lut_int_data : REG_lo_6;
  assign _0277_ = lo_wr_en_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6403" *) reg2dp_lut_int_data : REG_lo_5;
  assign _0266_ = lo_wr_en_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6341" *) reg2dp_lut_int_data : REG_lo_4;
  assign _0255_ = lo_wr_en_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6279" *) reg2dp_lut_int_data : REG_lo_3;
  assign _0244_ = lo_wr_en_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6217" *) reg2dp_lut_int_data : REG_lo_2;
  assign _0176_ = lo_wr_en_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6155" *) reg2dp_lut_int_data : REG_lo_1;
  assign _0065_ = lo_wr_en_0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:6093" *) reg2dp_lut_int_data : REG_lo_0;
  assign _0060_ = le_wr_en_64 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5839" *) reg2dp_lut_int_data : REG_le_64;
  assign _0059_ = le_wr_en_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5777" *) reg2dp_lut_int_data : REG_le_63;
  assign _0058_ = le_wr_en_62 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5715" *) reg2dp_lut_int_data : REG_le_62;
  assign _0057_ = le_wr_en_61 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5653" *) reg2dp_lut_int_data : REG_le_61;
  assign _0056_ = le_wr_en_60 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5591" *) reg2dp_lut_int_data : REG_le_60;
  assign _0054_ = le_wr_en_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5529" *) reg2dp_lut_int_data : REG_le_59;
  assign _0053_ = le_wr_en_58 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5467" *) reg2dp_lut_int_data : REG_le_58;
  assign _0052_ = le_wr_en_57 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5405" *) reg2dp_lut_int_data : REG_le_57;
  assign _0051_ = le_wr_en_56 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5343" *) reg2dp_lut_int_data : REG_le_56;
  assign _0050_ = le_wr_en_55 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5281" *) reg2dp_lut_int_data : REG_le_55;
  assign _0049_ = le_wr_en_54 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5219" *) reg2dp_lut_int_data : REG_le_54;
  assign _0048_ = le_wr_en_53 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5157" *) reg2dp_lut_int_data : REG_le_53;
  assign _0047_ = le_wr_en_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5095" *) reg2dp_lut_int_data : REG_le_52;
  assign _0046_ = le_wr_en_51 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:5033" *) reg2dp_lut_int_data : REG_le_51;
  assign _0045_ = le_wr_en_50 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4971" *) reg2dp_lut_int_data : REG_le_50;
  assign _0043_ = le_wr_en_49 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4909" *) reg2dp_lut_int_data : REG_le_49;
  assign _0042_ = le_wr_en_48 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4847" *) reg2dp_lut_int_data : REG_le_48;
  assign _0041_ = le_wr_en_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4785" *) reg2dp_lut_int_data : REG_le_47;
  assign _0040_ = le_wr_en_46 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4723" *) reg2dp_lut_int_data : REG_le_46;
  assign _0039_ = le_wr_en_45 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4661" *) reg2dp_lut_int_data : REG_le_45;
  assign _0038_ = le_wr_en_44 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4599" *) reg2dp_lut_int_data : REG_le_44;
  assign _0037_ = le_wr_en_43 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4537" *) reg2dp_lut_int_data : REG_le_43;
  assign _0036_ = le_wr_en_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4475" *) reg2dp_lut_int_data : REG_le_42;
  assign _0035_ = le_wr_en_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4413" *) reg2dp_lut_int_data : REG_le_41;
  assign _0034_ = le_wr_en_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4351" *) reg2dp_lut_int_data : REG_le_40;
  assign _0032_ = le_wr_en_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4289" *) reg2dp_lut_int_data : REG_le_39;
  assign _0031_ = le_wr_en_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4227" *) reg2dp_lut_int_data : REG_le_38;
  assign _0030_ = le_wr_en_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4165" *) reg2dp_lut_int_data : REG_le_37;
  assign _0029_ = le_wr_en_36 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4103" *) reg2dp_lut_int_data : REG_le_36;
  assign _0028_ = le_wr_en_35 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:4041" *) reg2dp_lut_int_data : REG_le_35;
  assign _0027_ = le_wr_en_34 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3979" *) reg2dp_lut_int_data : REG_le_34;
  assign _0026_ = le_wr_en_33 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3917" *) reg2dp_lut_int_data : REG_le_33;
  assign _0025_ = le_wr_en_32 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3855" *) reg2dp_lut_int_data : REG_le_32;
  assign _0024_ = le_wr_en_31 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3793" *) reg2dp_lut_int_data : REG_le_31;
  assign _0023_ = le_wr_en_30 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3731" *) reg2dp_lut_int_data : REG_le_30;
  assign _0021_ = le_wr_en_29 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3669" *) reg2dp_lut_int_data : REG_le_29;
  assign _0020_ = le_wr_en_28 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3607" *) reg2dp_lut_int_data : REG_le_28;
  assign _0019_ = le_wr_en_27 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3545" *) reg2dp_lut_int_data : REG_le_27;
  assign _0018_ = le_wr_en_26 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3483" *) reg2dp_lut_int_data : REG_le_26;
  assign _0017_ = le_wr_en_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3421" *) reg2dp_lut_int_data : REG_le_25;
  assign _0016_ = le_wr_en_24 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3359" *) reg2dp_lut_int_data : REG_le_24;
  assign _0015_ = le_wr_en_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3297" *) reg2dp_lut_int_data : REG_le_23;
  assign _0014_ = le_wr_en_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3235" *) reg2dp_lut_int_data : REG_le_22;
  assign _0013_ = le_wr_en_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3173" *) reg2dp_lut_int_data : REG_le_21;
  assign _0012_ = le_wr_en_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3111" *) reg2dp_lut_int_data : REG_le_20;
  assign _0010_ = le_wr_en_19 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:3049" *) reg2dp_lut_int_data : REG_le_19;
  assign _0009_ = le_wr_en_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2987" *) reg2dp_lut_int_data : REG_le_18;
  assign _0008_ = le_wr_en_17 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2925" *) reg2dp_lut_int_data : REG_le_17;
  assign _0007_ = le_wr_en_16 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2863" *) reg2dp_lut_int_data : REG_le_16;
  assign _0006_ = le_wr_en_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2801" *) reg2dp_lut_int_data : REG_le_15;
  assign _0005_ = le_wr_en_14 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2739" *) reg2dp_lut_int_data : REG_le_14;
  assign _0004_ = le_wr_en_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2677" *) reg2dp_lut_int_data : REG_le_13;
  assign _0003_ = le_wr_en_12 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2615" *) reg2dp_lut_int_data : REG_le_12;
  assign _0002_ = le_wr_en_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2553" *) reg2dp_lut_int_data : REG_le_11;
  assign _0001_ = le_wr_en_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2491" *) reg2dp_lut_int_data : REG_le_10;
  assign _0064_ = le_wr_en_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2429" *) reg2dp_lut_int_data : REG_le_9;
  assign _0063_ = le_wr_en_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2367" *) reg2dp_lut_int_data : REG_le_8;
  assign _0062_ = le_wr_en_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2305" *) reg2dp_lut_int_data : REG_le_7;
  assign _0061_ = le_wr_en_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2243" *) reg2dp_lut_int_data : REG_le_6;
  assign _0055_ = le_wr_en_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2181" *) reg2dp_lut_int_data : REG_le_5;
  assign _0044_ = le_wr_en_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2119" *) reg2dp_lut_int_data : REG_le_4;
  assign _0033_ = le_wr_en_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:2057" *) reg2dp_lut_int_data : REG_le_3;
  assign _0022_ = le_wr_en_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1995" *) reg2dp_lut_int_data : REG_le_2;
  assign _0011_ = le_wr_en_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1933" *) reg2dp_lut_int_data : REG_le_1;
  assign _0000_ = le_wr_en_0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1871" *) reg2dp_lut_int_data : REG_le_0;
  function [15:0] _6141_;
    input [15:0] a;
    input [4111:0] b;
    input [256:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1855|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1598" *)
    (* parallel_case *)
    casez (s)
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6141_ = b[15:0];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6141_ = b[31:16];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6141_ = b[47:32];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6141_ = b[63:48];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6141_ = b[79:64];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6141_ = b[95:80];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6141_ = b[111:96];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6141_ = b[127:112];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6141_ = b[143:128];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6141_ = b[159:144];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6141_ = b[175:160];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6141_ = b[191:176];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6141_ = b[207:192];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6141_ = b[223:208];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6141_ = b[239:224];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6141_ = b[255:240];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6141_ = b[271:256];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6141_ = b[287:272];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6141_ = b[303:288];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6141_ = b[319:304];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6141_ = b[335:320];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6141_ = b[351:336];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6141_ = b[367:352];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6141_ = b[383:368];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6141_ = b[399:384];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6141_ = b[415:400];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6141_ = b[431:416];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6141_ = b[447:432];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6141_ = b[463:448];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6141_ = b[479:464];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6141_ = b[495:480];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6141_ = b[511:496];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6141_ = b[527:512];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6141_ = b[543:528];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6141_ = b[559:544];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6141_ = b[575:560];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6141_ = b[591:576];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6141_ = b[607:592];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6141_ = b[623:608];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6141_ = b[639:624];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6141_ = b[655:640];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6141_ = b[671:656];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6141_ = b[687:672];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6141_ = b[703:688];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6141_ = b[719:704];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6141_ = b[735:720];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6141_ = b[751:736];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6141_ = b[767:752];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6141_ = b[783:768];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6141_ = b[799:784];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6141_ = b[815:800];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6141_ = b[831:816];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6141_ = b[847:832];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6141_ = b[863:848];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6141_ = b[879:864];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6141_ = b[895:880];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6141_ = b[911:896];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6141_ = b[927:912];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6141_ = b[943:928];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6141_ = b[959:944];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6141_ = b[975:960];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6141_ = b[991:976];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6141_ = b[1007:992];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6141_ = b[1023:1008];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6141_ = b[1039:1024];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6141_ = b[1055:1040];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6141_ = b[1071:1056];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6141_ = b[1087:1072];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6141_ = b[1103:1088];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6141_ = b[1119:1104];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6141_ = b[1135:1120];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6141_ = b[1151:1136];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1167:1152];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1183:1168];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1199:1184];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1215:1200];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1231:1216];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1247:1232];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1263:1248];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1279:1264];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1295:1280];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1311:1296];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1327:1312];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1343:1328];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1359:1344];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1375:1360];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1391:1376];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1407:1392];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1423:1408];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1439:1424];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1455:1440];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1471:1456];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1487:1472];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1503:1488];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1519:1504];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1535:1520];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1551:1536];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1567:1552];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1583:1568];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1599:1584];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1615:1600];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1631:1616];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1647:1632];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1663:1648];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1679:1664];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1695:1680];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1711:1696];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1727:1712];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1743:1728];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1759:1744];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1775:1760];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1791:1776];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1807:1792];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1823:1808];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1839:1824];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1855:1840];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1871:1856];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1887:1872];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1903:1888];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1919:1904];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1935:1920];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1951:1936];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1967:1952];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1983:1968];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[1999:1984];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2015:2000];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2031:2016];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2047:2032];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2063:2048];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2079:2064];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2095:2080];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2111:2096];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2127:2112];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2143:2128];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2159:2144];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2175:2160];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2191:2176];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2207:2192];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2223:2208];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2239:2224];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2255:2240];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2271:2256];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2287:2272];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2303:2288];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2319:2304];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2335:2320];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2351:2336];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2367:2352];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2383:2368];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2399:2384];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2415:2400];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2431:2416];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2447:2432];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2463:2448];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2479:2464];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2495:2480];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2511:2496];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2527:2512];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2543:2528];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2559:2544];
      257'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2575:2560];
      257'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2591:2576];
      257'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2607:2592];
      257'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2623:2608];
      257'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2639:2624];
      257'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2655:2640];
      257'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2671:2656];
      257'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2687:2672];
      257'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2703:2688];
      257'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2719:2704];
      257'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2735:2720];
      257'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2751:2736];
      257'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2767:2752];
      257'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2783:2768];
      257'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2799:2784];
      257'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2815:2800];
      257'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2831:2816];
      257'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2847:2832];
      257'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2863:2848];
      257'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2879:2864];
      257'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2895:2880];
      257'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2911:2896];
      257'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2927:2912];
      257'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2943:2928];
      257'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2959:2944];
      257'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2975:2960];
      257'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[2991:2976];
      257'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3007:2992];
      257'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3023:3008];
      257'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3039:3024];
      257'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3055:3040];
      257'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3071:3056];
      257'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3087:3072];
      257'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3103:3088];
      257'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3119:3104];
      257'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3135:3120];
      257'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3151:3136];
      257'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3167:3152];
      257'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3183:3168];
      257'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3199:3184];
      257'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3215:3200];
      257'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3231:3216];
      257'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3247:3232];
      257'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3263:3248];
      257'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3279:3264];
      257'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3295:3280];
      257'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3311:3296];
      257'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3327:3312];
      257'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3343:3328];
      257'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3359:3344];
      257'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3375:3360];
      257'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3391:3376];
      257'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3407:3392];
      257'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3423:3408];
      257'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3439:3424];
      257'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3455:3440];
      257'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3471:3456];
      257'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3487:3472];
      257'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3503:3488];
      257'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3519:3504];
      257'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3535:3520];
      257'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3551:3536];
      257'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3567:3552];
      257'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3583:3568];
      257'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3599:3584];
      257'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3615:3600];
      257'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3631:3616];
      257'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3647:3632];
      257'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3663:3648];
      257'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3679:3664];
      257'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3695:3680];
      257'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3711:3696];
      257'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3727:3712];
      257'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3743:3728];
      257'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3759:3744];
      257'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3775:3760];
      257'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3791:3776];
      257'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3807:3792];
      257'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3823:3808];
      257'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3839:3824];
      257'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3855:3840];
      257'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3871:3856];
      257'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3887:3872];
      257'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3903:3888];
      257'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3919:3904];
      257'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3935:3920];
      257'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3951:3936];
      257'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3967:3952];
      257'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3983:3968];
      257'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[3999:3984];
      257'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4015:4000];
      257'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4031:4016];
      257'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4047:4032];
      257'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4063:4048];
      257'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4079:4064];
      257'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4095:4080];
      257'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6141_ = b[4111:4096];
      default:
        _6141_ = a;
    endcase
  endfunction
  assign lo_lut_data = _6141_(16'b0000000000000000, { REG_lo_0, REG_lo_1, REG_lo_2, REG_lo_3, REG_lo_4, REG_lo_5, REG_lo_6, REG_lo_7, REG_lo_8, REG_lo_9, REG_lo_10, REG_lo_11, REG_lo_12, REG_lo_13, REG_lo_14, REG_lo_15, REG_lo_16, REG_lo_17, REG_lo_18, REG_lo_19, REG_lo_20, REG_lo_21, REG_lo_22, REG_lo_23, REG_lo_24, REG_lo_25, REG_lo_26, REG_lo_27, REG_lo_28, REG_lo_29, REG_lo_30, REG_lo_31, REG_lo_32, REG_lo_33, REG_lo_34, REG_lo_35, REG_lo_36, REG_lo_37, REG_lo_38, REG_lo_39, REG_lo_40, REG_lo_41, REG_lo_42, REG_lo_43, REG_lo_44, REG_lo_45, REG_lo_46, REG_lo_47, REG_lo_48, REG_lo_49, REG_lo_50, REG_lo_51, REG_lo_52, REG_lo_53, REG_lo_54, REG_lo_55, REG_lo_56, REG_lo_57, REG_lo_58, REG_lo_59, REG_lo_60, REG_lo_61, REG_lo_62, REG_lo_63, REG_lo_64, REG_lo_65, REG_lo_66, REG_lo_67, REG_lo_68, REG_lo_69, REG_lo_70, REG_lo_71, REG_lo_72, REG_lo_73, REG_lo_74, REG_lo_75, REG_lo_76, REG_lo_77, REG_lo_78, REG_lo_79, REG_lo_80, REG_lo_81, REG_lo_82, REG_lo_83, REG_lo_84, REG_lo_85, REG_lo_86, REG_lo_87, REG_lo_88, REG_lo_89, REG_lo_90, REG_lo_91, REG_lo_92, REG_lo_93, REG_lo_94, REG_lo_95, REG_lo_96, REG_lo_97, REG_lo_98, REG_lo_99, REG_lo_100, REG_lo_101, REG_lo_102, REG_lo_103, REG_lo_104, REG_lo_105, REG_lo_106, REG_lo_107, REG_lo_108, REG_lo_109, REG_lo_110, REG_lo_111, REG_lo_112, REG_lo_113, REG_lo_114, REG_lo_115, REG_lo_116, REG_lo_117, REG_lo_118, REG_lo_119, REG_lo_120, REG_lo_121, REG_lo_122, REG_lo_123, REG_lo_124, REG_lo_125, REG_lo_126, REG_lo_127, REG_lo_128, REG_lo_129, REG_lo_130, REG_lo_131, REG_lo_132, REG_lo_133, REG_lo_134, REG_lo_135, REG_lo_136, REG_lo_137, REG_lo_138, REG_lo_139, REG_lo_140, REG_lo_141, REG_lo_142, REG_lo_143, REG_lo_144, REG_lo_145, REG_lo_146, REG_lo_147, REG_lo_148, REG_lo_149, REG_lo_150, REG_lo_151, REG_lo_152, REG_lo_153, REG_lo_154, REG_lo_155, REG_lo_156, REG_lo_157, REG_lo_158, REG_lo_159, REG_lo_160, REG_lo_161, REG_lo_162, REG_lo_163, REG_lo_164, REG_lo_165, REG_lo_166, REG_lo_167, REG_lo_168, REG_lo_169, REG_lo_170, REG_lo_171, REG_lo_172, REG_lo_173, REG_lo_174, REG_lo_175, REG_lo_176, REG_lo_177, REG_lo_178, REG_lo_179, REG_lo_180, REG_lo_181, REG_lo_182, REG_lo_183, REG_lo_184, REG_lo_185, REG_lo_186, REG_lo_187, REG_lo_188, REG_lo_189, REG_lo_190, REG_lo_191, REG_lo_192, REG_lo_193, REG_lo_194, REG_lo_195, REG_lo_196, REG_lo_197, REG_lo_198, REG_lo_199, REG_lo_200, REG_lo_201, REG_lo_202, REG_lo_203, REG_lo_204, REG_lo_205, REG_lo_206, REG_lo_207, REG_lo_208, REG_lo_209, REG_lo_210, REG_lo_211, REG_lo_212, REG_lo_213, REG_lo_214, REG_lo_215, REG_lo_216, REG_lo_217, REG_lo_218, REG_lo_219, REG_lo_220, REG_lo_221, REG_lo_222, REG_lo_223, REG_lo_224, REG_lo_225, REG_lo_226, REG_lo_227, REG_lo_228, REG_lo_229, REG_lo_230, REG_lo_231, REG_lo_232, REG_lo_233, REG_lo_234, REG_lo_235, REG_lo_236, REG_lo_237, REG_lo_238, REG_lo_239, REG_lo_240, REG_lo_241, REG_lo_242, REG_lo_243, REG_lo_244, REG_lo_245, REG_lo_246, REG_lo_247, REG_lo_248, REG_lo_249, REG_lo_250, REG_lo_251, REG_lo_252, REG_lo_253, REG_lo_254, REG_lo_255, REG_lo_256 }, { _0527_, _0538_, _0549_, _0560_, _0571_, _0582_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0603_, _0604_, _0605_, _0606_, _0607_, _0608_, _0609_, _0610_, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0388_, _0389_, _0390_, _0391_, _0392_, _0393_, _0394_, _0395_, _0396_, _0397_, _0398_, _0399_, _0400_, _0401_, _0402_, _0403_, _0404_, _0405_, _0406_, _0407_, _0408_, _0409_, _0410_, _0411_, _0412_, _0413_, _0414_, _0415_, _0416_, _0417_, _0418_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_, _0451_, _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0484_, _0485_, _0486_, _0487_, _0488_, _0489_, _0490_, _0491_, _0492_, _0493_, _0494_, _0495_, _0496_, _0497_, _0498_, _0499_, _0500_, _0501_, _0502_, _0503_, _0504_, _0505_, _0506_, _0507_, _0508_, _0509_, _0510_, _0511_, _0512_, _0513_, _0514_, _0515_, _0516_, _0517_, _0518_, _0519_, _0520_, _0521_, _0522_, _0523_, _0524_, _0525_, _0526_, _0528_, _0529_, _0530_, _0531_, _0532_, _0533_, _0534_, _0535_, _0536_, _0537_, _0539_, _0540_, _0541_, _0542_, _0543_, _0544_, _0545_, _0546_, _0547_, _0548_, _0550_, _0551_, _0552_, _0553_, _0554_, _0555_, _0556_, _0557_, _0558_, _0559_, _0561_, _0562_, _0563_, _0564_, _0565_, _0566_, _0567_, _0568_, _0569_, _0570_, _0572_, _0573_, _0574_, _0575_, _0576_, _0577_, _0578_, _0579_, _0580_, _0581_, _0583_, _0584_, _0585_, _0586_ });
  function [15:0] _6142_;
    input [15:0] a;
    input [1039:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1330|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1265" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _6142_ = b[15:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _6142_ = b[31:16];
      65'b??????????????????????????????????????????????????????????????1??:
        _6142_ = b[47:32];
      65'b?????????????????????????????????????????????????????????????1???:
        _6142_ = b[63:48];
      65'b????????????????????????????????????????????????????????????1????:
        _6142_ = b[79:64];
      65'b???????????????????????????????????????????????????????????1?????:
        _6142_ = b[95:80];
      65'b??????????????????????????????????????????????????????????1??????:
        _6142_ = b[111:96];
      65'b?????????????????????????????????????????????????????????1???????:
        _6142_ = b[127:112];
      65'b????????????????????????????????????????????????????????1????????:
        _6142_ = b[143:128];
      65'b???????????????????????????????????????????????????????1?????????:
        _6142_ = b[159:144];
      65'b??????????????????????????????????????????????????????1??????????:
        _6142_ = b[175:160];
      65'b?????????????????????????????????????????????????????1???????????:
        _6142_ = b[191:176];
      65'b????????????????????????????????????????????????????1????????????:
        _6142_ = b[207:192];
      65'b???????????????????????????????????????????????????1?????????????:
        _6142_ = b[223:208];
      65'b??????????????????????????????????????????????????1??????????????:
        _6142_ = b[239:224];
      65'b?????????????????????????????????????????????????1???????????????:
        _6142_ = b[255:240];
      65'b????????????????????????????????????????????????1????????????????:
        _6142_ = b[271:256];
      65'b???????????????????????????????????????????????1?????????????????:
        _6142_ = b[287:272];
      65'b??????????????????????????????????????????????1??????????????????:
        _6142_ = b[303:288];
      65'b?????????????????????????????????????????????1???????????????????:
        _6142_ = b[319:304];
      65'b????????????????????????????????????????????1????????????????????:
        _6142_ = b[335:320];
      65'b???????????????????????????????????????????1?????????????????????:
        _6142_ = b[351:336];
      65'b??????????????????????????????????????????1??????????????????????:
        _6142_ = b[367:352];
      65'b?????????????????????????????????????????1???????????????????????:
        _6142_ = b[383:368];
      65'b????????????????????????????????????????1????????????????????????:
        _6142_ = b[399:384];
      65'b???????????????????????????????????????1?????????????????????????:
        _6142_ = b[415:400];
      65'b??????????????????????????????????????1??????????????????????????:
        _6142_ = b[431:416];
      65'b?????????????????????????????????????1???????????????????????????:
        _6142_ = b[447:432];
      65'b????????????????????????????????????1????????????????????????????:
        _6142_ = b[463:448];
      65'b???????????????????????????????????1?????????????????????????????:
        _6142_ = b[479:464];
      65'b??????????????????????????????????1??????????????????????????????:
        _6142_ = b[495:480];
      65'b?????????????????????????????????1???????????????????????????????:
        _6142_ = b[511:496];
      65'b????????????????????????????????1????????????????????????????????:
        _6142_ = b[527:512];
      65'b???????????????????????????????1?????????????????????????????????:
        _6142_ = b[543:528];
      65'b??????????????????????????????1??????????????????????????????????:
        _6142_ = b[559:544];
      65'b?????????????????????????????1???????????????????????????????????:
        _6142_ = b[575:560];
      65'b????????????????????????????1????????????????????????????????????:
        _6142_ = b[591:576];
      65'b???????????????????????????1?????????????????????????????????????:
        _6142_ = b[607:592];
      65'b??????????????????????????1??????????????????????????????????????:
        _6142_ = b[623:608];
      65'b?????????????????????????1???????????????????????????????????????:
        _6142_ = b[639:624];
      65'b????????????????????????1????????????????????????????????????????:
        _6142_ = b[655:640];
      65'b???????????????????????1?????????????????????????????????????????:
        _6142_ = b[671:656];
      65'b??????????????????????1??????????????????????????????????????????:
        _6142_ = b[687:672];
      65'b?????????????????????1???????????????????????????????????????????:
        _6142_ = b[703:688];
      65'b????????????????????1????????????????????????????????????????????:
        _6142_ = b[719:704];
      65'b???????????????????1?????????????????????????????????????????????:
        _6142_ = b[735:720];
      65'b??????????????????1??????????????????????????????????????????????:
        _6142_ = b[751:736];
      65'b?????????????????1???????????????????????????????????????????????:
        _6142_ = b[767:752];
      65'b????????????????1????????????????????????????????????????????????:
        _6142_ = b[783:768];
      65'b???????????????1?????????????????????????????????????????????????:
        _6142_ = b[799:784];
      65'b??????????????1??????????????????????????????????????????????????:
        _6142_ = b[815:800];
      65'b?????????????1???????????????????????????????????????????????????:
        _6142_ = b[831:816];
      65'b????????????1????????????????????????????????????????????????????:
        _6142_ = b[847:832];
      65'b???????????1?????????????????????????????????????????????????????:
        _6142_ = b[863:848];
      65'b??????????1??????????????????????????????????????????????????????:
        _6142_ = b[879:864];
      65'b?????????1???????????????????????????????????????????????????????:
        _6142_ = b[895:880];
      65'b????????1????????????????????????????????????????????????????????:
        _6142_ = b[911:896];
      65'b???????1?????????????????????????????????????????????????????????:
        _6142_ = b[927:912];
      65'b??????1??????????????????????????????????????????????????????????:
        _6142_ = b[943:928];
      65'b?????1???????????????????????????????????????????????????????????:
        _6142_ = b[959:944];
      65'b????1????????????????????????????????????????????????????????????:
        _6142_ = b[975:960];
      65'b???1?????????????????????????????????????????????????????????????:
        _6142_ = b[991:976];
      65'b??1??????????????????????????????????????????????????????????????:
        _6142_ = b[1007:992];
      65'b?1???????????????????????????????????????????????????????????????:
        _6142_ = b[1023:1008];
      65'b1????????????????????????????????????????????????????????????????:
        _6142_ = b[1039:1024];
      default:
        _6142_ = a;
    endcase
  endfunction
  assign le_lut_data = _6142_(16'b0000000000000000, { REG_le_0, REG_le_1, REG_le_2, REG_le_3, REG_le_4, REG_le_5, REG_le_6, REG_le_7, REG_le_8, REG_le_9, REG_le_10, REG_le_11, REG_le_12, REG_le_13, REG_le_14, REG_le_15, REG_le_16, REG_le_17, REG_le_18, REG_le_19, REG_le_20, REG_le_21, REG_le_22, REG_le_23, REG_le_24, REG_le_25, REG_le_26, REG_le_27, REG_le_28, REG_le_29, REG_le_30, REG_le_31, REG_le_32, REG_le_33, REG_le_34, REG_le_35, REG_le_36, REG_le_37, REG_le_38, REG_le_39, REG_le_40, REG_le_41, REG_le_42, REG_le_43, REG_le_44, REG_le_45, REG_le_46, REG_le_47, REG_le_48, REG_le_49, REG_le_50, REG_le_51, REG_le_52, REG_le_53, REG_le_54, REG_le_55, REG_le_56, REG_le_57, REG_le_58, REG_le_59, REG_le_60, REG_le_61, REG_le_62, REG_le_63, REG_le_64 }, { _0527_, _0538_, _0549_, _0560_, _0571_, _0582_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0603_, _0604_, _0605_, _0606_, _0607_, _0608_, _0609_, _0610_, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0388_ });
  assign _2709_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22381" *) { perf_lut_oflow_cnt_cur[0], perf_lut_oflow_cnt_cur[1], perf_lut_oflow_cnt_cur[2], perf_lut_oflow_cnt_cur[3], perf_lut_oflow_cnt_cur[4], perf_lut_oflow_cnt_cur[5], perf_lut_oflow_cnt_cur[6], perf_lut_oflow_cnt_cur[7], perf_lut_oflow_cnt_cur[8], perf_lut_oflow_cnt_cur[9], perf_lut_oflow_cnt_cur[10], perf_lut_oflow_cnt_cur[11], perf_lut_oflow_cnt_cur[12], perf_lut_oflow_cnt_cur[13], perf_lut_oflow_cnt_cur[14], perf_lut_oflow_cnt_cur[15], perf_lut_oflow_cnt_cur[16], perf_lut_oflow_cnt_cur[17], perf_lut_oflow_cnt_cur[18], perf_lut_oflow_cnt_cur[19], perf_lut_oflow_cnt_cur[20], perf_lut_oflow_cnt_cur[21], perf_lut_oflow_cnt_cur[22], perf_lut_oflow_cnt_cur[23], perf_lut_oflow_cnt_cur[24], perf_lut_oflow_cnt_cur[25], perf_lut_oflow_cnt_cur[26], perf_lut_oflow_cnt_cur[27], perf_lut_oflow_cnt_cur[28], perf_lut_oflow_cnt_cur[29], perf_lut_oflow_cnt_cur[30], perf_lut_oflow_cnt_cur[31] };
  assign _2710_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22424" *) { perf_lut_uflow_cnt_cur[0], perf_lut_uflow_cnt_cur[1], perf_lut_uflow_cnt_cur[2], perf_lut_uflow_cnt_cur[3], perf_lut_uflow_cnt_cur[4], perf_lut_uflow_cnt_cur[5], perf_lut_uflow_cnt_cur[6], perf_lut_uflow_cnt_cur[7], perf_lut_uflow_cnt_cur[8], perf_lut_uflow_cnt_cur[9], perf_lut_uflow_cnt_cur[10], perf_lut_uflow_cnt_cur[11], perf_lut_uflow_cnt_cur[12], perf_lut_uflow_cnt_cur[13], perf_lut_uflow_cnt_cur[14], perf_lut_uflow_cnt_cur[15], perf_lut_uflow_cnt_cur[16], perf_lut_uflow_cnt_cur[17], perf_lut_uflow_cnt_cur[18], perf_lut_uflow_cnt_cur[19], perf_lut_uflow_cnt_cur[20], perf_lut_uflow_cnt_cur[21], perf_lut_uflow_cnt_cur[22], perf_lut_uflow_cnt_cur[23], perf_lut_uflow_cnt_cur[24], perf_lut_uflow_cnt_cur[25], perf_lut_uflow_cnt_cur[26], perf_lut_uflow_cnt_cur[27], perf_lut_uflow_cnt_cur[28], perf_lut_uflow_cnt_cur[29], perf_lut_uflow_cnt_cur[30], perf_lut_uflow_cnt_cur[31] };
  assign _2711_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22471" *) { perf_lut_hybrid_cnt_cur[0], perf_lut_hybrid_cnt_cur[1], perf_lut_hybrid_cnt_cur[2], perf_lut_hybrid_cnt_cur[3], perf_lut_hybrid_cnt_cur[4], perf_lut_hybrid_cnt_cur[5], perf_lut_hybrid_cnt_cur[6], perf_lut_hybrid_cnt_cur[7], perf_lut_hybrid_cnt_cur[8], perf_lut_hybrid_cnt_cur[9], perf_lut_hybrid_cnt_cur[10], perf_lut_hybrid_cnt_cur[11], perf_lut_hybrid_cnt_cur[12], perf_lut_hybrid_cnt_cur[13], perf_lut_hybrid_cnt_cur[14], perf_lut_hybrid_cnt_cur[15], perf_lut_hybrid_cnt_cur[16], perf_lut_hybrid_cnt_cur[17], perf_lut_hybrid_cnt_cur[18], perf_lut_hybrid_cnt_cur[19], perf_lut_hybrid_cnt_cur[20], perf_lut_hybrid_cnt_cur[21], perf_lut_hybrid_cnt_cur[22], perf_lut_hybrid_cnt_cur[23], perf_lut_hybrid_cnt_cur[24], perf_lut_hybrid_cnt_cur[25], perf_lut_hybrid_cnt_cur[26], perf_lut_hybrid_cnt_cur[27], perf_lut_hybrid_cnt_cur[28], perf_lut_hybrid_cnt_cur[29], perf_lut_hybrid_cnt_cur[30], perf_lut_hybrid_cnt_cur[31] };
  assign _2712_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22514" *) { perf_lut_le_hit_cnt_cur[0], perf_lut_le_hit_cnt_cur[1], perf_lut_le_hit_cnt_cur[2], perf_lut_le_hit_cnt_cur[3], perf_lut_le_hit_cnt_cur[4], perf_lut_le_hit_cnt_cur[5], perf_lut_le_hit_cnt_cur[6], perf_lut_le_hit_cnt_cur[7], perf_lut_le_hit_cnt_cur[8], perf_lut_le_hit_cnt_cur[9], perf_lut_le_hit_cnt_cur[10], perf_lut_le_hit_cnt_cur[11], perf_lut_le_hit_cnt_cur[12], perf_lut_le_hit_cnt_cur[13], perf_lut_le_hit_cnt_cur[14], perf_lut_le_hit_cnt_cur[15], perf_lut_le_hit_cnt_cur[16], perf_lut_le_hit_cnt_cur[17], perf_lut_le_hit_cnt_cur[18], perf_lut_le_hit_cnt_cur[19], perf_lut_le_hit_cnt_cur[20], perf_lut_le_hit_cnt_cur[21], perf_lut_le_hit_cnt_cur[22], perf_lut_le_hit_cnt_cur[23], perf_lut_le_hit_cnt_cur[24], perf_lut_le_hit_cnt_cur[25], perf_lut_le_hit_cnt_cur[26], perf_lut_le_hit_cnt_cur[27], perf_lut_le_hit_cnt_cur[28], perf_lut_le_hit_cnt_cur[29], perf_lut_le_hit_cnt_cur[30], perf_lut_le_hit_cnt_cur[31] };
  assign _2713_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22557" *) { perf_lut_lo_hit_cnt_cur[0], perf_lut_lo_hit_cnt_cur[1], perf_lut_lo_hit_cnt_cur[2], perf_lut_lo_hit_cnt_cur[3], perf_lut_lo_hit_cnt_cur[4], perf_lut_lo_hit_cnt_cur[5], perf_lut_lo_hit_cnt_cur[6], perf_lut_lo_hit_cnt_cur[7], perf_lut_lo_hit_cnt_cur[8], perf_lut_lo_hit_cnt_cur[9], perf_lut_lo_hit_cnt_cur[10], perf_lut_lo_hit_cnt_cur[11], perf_lut_lo_hit_cnt_cur[12], perf_lut_lo_hit_cnt_cur[13], perf_lut_lo_hit_cnt_cur[14], perf_lut_lo_hit_cnt_cur[15], perf_lut_lo_hit_cnt_cur[16], perf_lut_lo_hit_cnt_cur[17], perf_lut_lo_hit_cnt_cur[18], perf_lut_lo_hit_cnt_cur[19], perf_lut_lo_hit_cnt_cur[20], perf_lut_lo_hit_cnt_cur[21], perf_lut_lo_hit_cnt_cur[22], perf_lut_lo_hit_cnt_cur[23], perf_lut_lo_hit_cnt_cur[24], perf_lut_lo_hit_cnt_cur[25], perf_lut_lo_hit_cnt_cur[26], perf_lut_lo_hit_cnt_cur[27], perf_lut_lo_hit_cnt_cur[28], perf_lut_lo_hit_cnt_cur[29], perf_lut_lo_hit_cnt_cur[30], perf_lut_lo_hit_cnt_cur[31] };
  assign _2714_ = $signed(2'b01) << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31132" *) reg2dp_lut_le_index_offset;
  assign dp2reg_lut_int_data = reg2dp_lut_int_table_id ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:1863" *) lo_lut_data : le_lut_data;
  assign _0324_ = p1_pipe_ready_bc ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22225" *) idx2lut_pvld : 1'b1;
  assign _0323_ = _0646_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22230" *) idx2lut_pd : p1_pipe_data;
  assign perf_lut_oflow_add = _2709_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22381" *) 3'b000 : lut_oflow_sum;
  assign perf_lut_oflow_cnt_new = perf_lut_oflow_adv ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22402" *) perf_lut_oflow_cnt_mod : perf_lut_oflow_cnt_cur;
  assign perf_lut_oflow_cnt_nxt = op_en_load ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22403" *) 32'd0 : perf_lut_oflow_cnt_new;
  assign perf_lut_uflow_add = _2710_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22424" *) 3'b000 : lut_uflow_sum;
  assign perf_lut_uflow_cnt_new = perf_lut_uflow_adv ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22445" *) perf_lut_uflow_cnt_mod : perf_lut_uflow_cnt_cur;
  assign perf_lut_uflow_cnt_nxt = op_en_load ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22446" *) 32'd0 : perf_lut_uflow_cnt_new;
  assign perf_lut_hybrid_add = _2711_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22471" *) 3'b000 : lut_hybrid_sum;
  assign perf_lut_hybrid_cnt_new = perf_lut_hybrid_adv ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22492" *) perf_lut_hybrid_cnt_mod : perf_lut_hybrid_cnt_cur;
  assign perf_lut_hybrid_cnt_nxt = op_en_load ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22493" *) 32'd0 : perf_lut_hybrid_cnt_new;
  assign perf_lut_le_hit_add = _2712_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22514" *) 3'b000 : lut_le_hit_sum;
  assign perf_lut_le_hit_cnt_new = perf_lut_le_hit_adv ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22535" *) perf_lut_le_hit_cnt_mod : perf_lut_le_hit_cnt_cur;
  assign perf_lut_le_hit_cnt_nxt = op_en_load ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22536" *) 32'd0 : perf_lut_le_hit_cnt_new;
  assign perf_lut_lo_hit_add = _2713_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22557" *) 3'b000 : lut_lo_hit_sum;
  assign perf_lut_lo_hit_cnt_new = perf_lut_lo_hit_adv ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22578" *) perf_lut_lo_hit_cnt_mod : perf_lut_lo_hit_cnt_cur;
  assign perf_lut_lo_hit_cnt_nxt = op_en_load ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:22579" *) 32'd0 : perf_lut_lo_hit_cnt_new;
  assign dat_in_y0_0 = p1_pipe_data[276] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30992" *) lo_data0_0 : le_data0_0;
  assign dat_in_y0_1 = p1_pipe_data[277] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30993" *) lo_data0_1 : le_data0_1;
  assign dat_in_y0_2 = p1_pipe_data[278] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30994" *) lo_data0_2 : le_data0_2;
  assign dat_in_y0_3 = p1_pipe_data[279] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30995" *) lo_data0_3 : le_data0_3;
  assign dat_in_y1_0 = p1_pipe_data[276] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30996" *) lo_data1_0 : le_data1_0;
  assign dat_in_y1_1 = p1_pipe_data[277] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30997" *) lo_data1_1 : le_data1_1;
  assign dat_in_y1_2 = p1_pipe_data[278] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30998" *) lo_data1_2 : le_data1_2;
  assign dat_in_y1_3 = p1_pipe_data[279] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:30999" *) lo_data1_3 : le_data1_3;
  assign _2715_ = reg2dp_lut_le_index_offset[7] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31132" *) 32'd0 : _2714_;
  assign _0326_ = dat_fifo_rd_prdy ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31589" *) dat_fifo_rd_pvld : 1'b1;
  assign _0325_ = _0647_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31594" *) { out_flow3, out_flow2, out_flow1, out_flow0, out_bias3, out_bias2, out_bias1, out_bias0, out_offset3, out_offset2, out_offset1, out_offset0, out_shift3, out_shift2, out_shift1, out_shift0, out_scale3, out_scale2, out_scale1, out_scale0, dat_fifo_rd_pd, cmd_fifo_rd_pd[139:0], cmd_fifo_rd_pd[267:140] } : p2_pipe_data;
  assign p2_skid_ready = p2_skid_valid ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31610" *) lut2inp_prdy : _0652_;
  assign _0328_ = p2_skid_valid ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31618" *) _0651_ : p2_skid_catch;
  assign _0327_ = p2_skid_catch ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31625" *) p2_pipe_data : p2_skid_data;
  assign lut2inp_pvld = p2_pipe_ready ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31635" *) p2_pipe_valid : p2_skid_valid;
  assign lut2inp_pd = p2_pipe_ready ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31637" *) p2_pipe_data : p2_skid_data;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31051" *)
  NV_NVDLA_SDP_CORE_Y_LUT_cmd u_cmd (
    .cmd_fifo_rd_pd(cmd_fifo_rd_pd),
    .cmd_fifo_rd_prdy(cmd_fifo_rd_prdy),
    .cmd_fifo_rd_pvld(cmd_fifo_rd_pvld),
    .cmd_fifo_wr_pd(p1_pipe_data[279:0]),
    .cmd_fifo_wr_prdy(cmd_fifo_wr_prdy),
    .cmd_fifo_wr_pvld(p1_pipe_valid),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn),
    .pwrbus_ram_pd(pwrbus_ram_pd)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_lut.v:31013" *)
  NV_NVDLA_SDP_CORE_Y_LUT_dat u_dat (
    .dat_fifo_rd_pd(dat_fifo_rd_pd),
    .dat_fifo_rd_prdy(dat_fifo_rd_prdy),
    .dat_fifo_rd_pvld(dat_fifo_rd_pvld),
    .dat_fifo_wr_pd({ dat_in_y1_3, dat_in_y1_2, dat_in_y1_1, dat_in_y1_0, dat_in_y0_3, dat_in_y0_2, dat_in_y0_1, dat_in_y0_0 }),
    .dat_fifo_wr_pvld(dat_fifo_wr_pvld),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn),
    .pwrbus_ram_pd(pwrbus_ram_pd)
  );
  assign REG_le_100 = 16'b0000000000000000;
  assign REG_le_101 = 16'b0000000000000000;
  assign REG_le_102 = 16'b0000000000000000;
  assign REG_le_103 = 16'b0000000000000000;
  assign REG_le_104 = 16'b0000000000000000;
  assign REG_le_105 = 16'b0000000000000000;
  assign REG_le_106 = 16'b0000000000000000;
  assign REG_le_107 = 16'b0000000000000000;
  assign REG_le_108 = 16'b0000000000000000;
  assign REG_le_109 = 16'b0000000000000000;
  assign REG_le_110 = 16'b0000000000000000;
  assign REG_le_111 = 16'b0000000000000000;
  assign REG_le_112 = 16'b0000000000000000;
  assign REG_le_113 = 16'b0000000000000000;
  assign REG_le_114 = 16'b0000000000000000;
  assign REG_le_115 = 16'b0000000000000000;
  assign REG_le_116 = 16'b0000000000000000;
  assign REG_le_117 = 16'b0000000000000000;
  assign REG_le_118 = 16'b0000000000000000;
  assign REG_le_119 = 16'b0000000000000000;
  assign REG_le_120 = 16'b0000000000000000;
  assign REG_le_121 = 16'b0000000000000000;
  assign REG_le_122 = 16'b0000000000000000;
  assign REG_le_123 = 16'b0000000000000000;
  assign REG_le_124 = 16'b0000000000000000;
  assign REG_le_125 = 16'b0000000000000000;
  assign REG_le_126 = 16'b0000000000000000;
  assign REG_le_127 = 16'b0000000000000000;
  assign REG_le_128 = 16'b0000000000000000;
  assign REG_le_129 = 16'b0000000000000000;
  assign REG_le_130 = 16'b0000000000000000;
  assign REG_le_131 = 16'b0000000000000000;
  assign REG_le_132 = 16'b0000000000000000;
  assign REG_le_133 = 16'b0000000000000000;
  assign REG_le_134 = 16'b0000000000000000;
  assign REG_le_135 = 16'b0000000000000000;
  assign REG_le_136 = 16'b0000000000000000;
  assign REG_le_137 = 16'b0000000000000000;
  assign REG_le_138 = 16'b0000000000000000;
  assign REG_le_139 = 16'b0000000000000000;
  assign REG_le_140 = 16'b0000000000000000;
  assign REG_le_141 = 16'b0000000000000000;
  assign REG_le_142 = 16'b0000000000000000;
  assign REG_le_143 = 16'b0000000000000000;
  assign REG_le_144 = 16'b0000000000000000;
  assign REG_le_145 = 16'b0000000000000000;
  assign REG_le_146 = 16'b0000000000000000;
  assign REG_le_147 = 16'b0000000000000000;
  assign REG_le_148 = 16'b0000000000000000;
  assign REG_le_149 = 16'b0000000000000000;
  assign REG_le_150 = 16'b0000000000000000;
  assign REG_le_151 = 16'b0000000000000000;
  assign REG_le_152 = 16'b0000000000000000;
  assign REG_le_153 = 16'b0000000000000000;
  assign REG_le_154 = 16'b0000000000000000;
  assign REG_le_155 = 16'b0000000000000000;
  assign REG_le_156 = 16'b0000000000000000;
  assign REG_le_157 = 16'b0000000000000000;
  assign REG_le_158 = 16'b0000000000000000;
  assign REG_le_159 = 16'b0000000000000000;
  assign REG_le_160 = 16'b0000000000000000;
  assign REG_le_161 = 16'b0000000000000000;
  assign REG_le_162 = 16'b0000000000000000;
  assign REG_le_163 = 16'b0000000000000000;
  assign REG_le_164 = 16'b0000000000000000;
  assign REG_le_165 = 16'b0000000000000000;
  assign REG_le_166 = 16'b0000000000000000;
  assign REG_le_167 = 16'b0000000000000000;
  assign REG_le_168 = 16'b0000000000000000;
  assign REG_le_169 = 16'b0000000000000000;
  assign REG_le_170 = 16'b0000000000000000;
  assign REG_le_171 = 16'b0000000000000000;
  assign REG_le_172 = 16'b0000000000000000;
  assign REG_le_173 = 16'b0000000000000000;
  assign REG_le_174 = 16'b0000000000000000;
  assign REG_le_175 = 16'b0000000000000000;
  assign REG_le_176 = 16'b0000000000000000;
  assign REG_le_177 = 16'b0000000000000000;
  assign REG_le_178 = 16'b0000000000000000;
  assign REG_le_179 = 16'b0000000000000000;
  assign REG_le_180 = 16'b0000000000000000;
  assign REG_le_181 = 16'b0000000000000000;
  assign REG_le_182 = 16'b0000000000000000;
  assign REG_le_183 = 16'b0000000000000000;
  assign REG_le_184 = 16'b0000000000000000;
  assign REG_le_185 = 16'b0000000000000000;
  assign REG_le_186 = 16'b0000000000000000;
  assign REG_le_187 = 16'b0000000000000000;
  assign REG_le_188 = 16'b0000000000000000;
  assign REG_le_189 = 16'b0000000000000000;
  assign REG_le_190 = 16'b0000000000000000;
  assign REG_le_191 = 16'b0000000000000000;
  assign REG_le_192 = 16'b0000000000000000;
  assign REG_le_193 = 16'b0000000000000000;
  assign REG_le_194 = 16'b0000000000000000;
  assign REG_le_195 = 16'b0000000000000000;
  assign REG_le_196 = 16'b0000000000000000;
  assign REG_le_197 = 16'b0000000000000000;
  assign REG_le_198 = 16'b0000000000000000;
  assign REG_le_199 = 16'b0000000000000000;
  assign REG_le_200 = 16'b0000000000000000;
  assign REG_le_201 = 16'b0000000000000000;
  assign REG_le_202 = 16'b0000000000000000;
  assign REG_le_203 = 16'b0000000000000000;
  assign REG_le_204 = 16'b0000000000000000;
  assign REG_le_205 = 16'b0000000000000000;
  assign REG_le_206 = 16'b0000000000000000;
  assign REG_le_207 = 16'b0000000000000000;
  assign REG_le_208 = 16'b0000000000000000;
  assign REG_le_209 = 16'b0000000000000000;
  assign REG_le_210 = 16'b0000000000000000;
  assign REG_le_211 = 16'b0000000000000000;
  assign REG_le_212 = 16'b0000000000000000;
  assign REG_le_213 = 16'b0000000000000000;
  assign REG_le_214 = 16'b0000000000000000;
  assign REG_le_215 = 16'b0000000000000000;
  assign REG_le_216 = 16'b0000000000000000;
  assign REG_le_217 = 16'b0000000000000000;
  assign REG_le_218 = 16'b0000000000000000;
  assign REG_le_219 = 16'b0000000000000000;
  assign REG_le_220 = 16'b0000000000000000;
  assign REG_le_221 = 16'b0000000000000000;
  assign REG_le_222 = 16'b0000000000000000;
  assign REG_le_223 = 16'b0000000000000000;
  assign REG_le_224 = 16'b0000000000000000;
  assign REG_le_225 = 16'b0000000000000000;
  assign REG_le_226 = 16'b0000000000000000;
  assign REG_le_227 = 16'b0000000000000000;
  assign REG_le_228 = 16'b0000000000000000;
  assign REG_le_229 = 16'b0000000000000000;
  assign REG_le_230 = 16'b0000000000000000;
  assign REG_le_231 = 16'b0000000000000000;
  assign REG_le_232 = 16'b0000000000000000;
  assign REG_le_233 = 16'b0000000000000000;
  assign REG_le_234 = 16'b0000000000000000;
  assign REG_le_235 = 16'b0000000000000000;
  assign REG_le_236 = 16'b0000000000000000;
  assign REG_le_237 = 16'b0000000000000000;
  assign REG_le_238 = 16'b0000000000000000;
  assign REG_le_239 = 16'b0000000000000000;
  assign REG_le_240 = 16'b0000000000000000;
  assign REG_le_241 = 16'b0000000000000000;
  assign REG_le_242 = 16'b0000000000000000;
  assign REG_le_243 = 16'b0000000000000000;
  assign REG_le_244 = 16'b0000000000000000;
  assign REG_le_245 = 16'b0000000000000000;
  assign REG_le_246 = 16'b0000000000000000;
  assign REG_le_247 = 16'b0000000000000000;
  assign REG_le_248 = 16'b0000000000000000;
  assign REG_le_249 = 16'b0000000000000000;
  assign REG_le_250 = 16'b0000000000000000;
  assign REG_le_251 = 16'b0000000000000000;
  assign REG_le_252 = 16'b0000000000000000;
  assign REG_le_253 = 16'b0000000000000000;
  assign REG_le_254 = 16'b0000000000000000;
  assign REG_le_255 = 16'b0000000000000000;
  assign REG_le_256 = 16'b0000000000000000;
  assign REG_le_65 = 16'b0000000000000000;
  assign REG_le_66 = 16'b0000000000000000;
  assign REG_le_67 = 16'b0000000000000000;
  assign REG_le_68 = 16'b0000000000000000;
  assign REG_le_69 = 16'b0000000000000000;
  assign REG_le_70 = 16'b0000000000000000;
  assign REG_le_71 = 16'b0000000000000000;
  assign REG_le_72 = 16'b0000000000000000;
  assign REG_le_73 = 16'b0000000000000000;
  assign REG_le_74 = 16'b0000000000000000;
  assign REG_le_75 = 16'b0000000000000000;
  assign REG_le_76 = 16'b0000000000000000;
  assign REG_le_77 = 16'b0000000000000000;
  assign REG_le_78 = 16'b0000000000000000;
  assign REG_le_79 = 16'b0000000000000000;
  assign REG_le_80 = 16'b0000000000000000;
  assign REG_le_81 = 16'b0000000000000000;
  assign REG_le_82 = 16'b0000000000000000;
  assign REG_le_83 = 16'b0000000000000000;
  assign REG_le_84 = 16'b0000000000000000;
  assign REG_le_85 = 16'b0000000000000000;
  assign REG_le_86 = 16'b0000000000000000;
  assign REG_le_87 = 16'b0000000000000000;
  assign REG_le_88 = 16'b0000000000000000;
  assign REG_le_89 = 16'b0000000000000000;
  assign REG_le_90 = 16'b0000000000000000;
  assign REG_le_91 = 16'b0000000000000000;
  assign REG_le_92 = 16'b0000000000000000;
  assign REG_le_93 = 16'b0000000000000000;
  assign REG_le_94 = 16'b0000000000000000;
  assign REG_le_95 = 16'b0000000000000000;
  assign REG_le_96 = 16'b0000000000000000;
  assign REG_le_97 = 16'b0000000000000000;
  assign REG_le_98 = 16'b0000000000000000;
  assign REG_le_99 = 16'b0000000000000000;
  assign cmd_fifo_wr_pd = p1_pipe_data[279:0];
  assign cmd_fifo_wr_pvld = p1_pipe_valid;
  assign dat_fifo_wr_pd = { dat_in_y1_3, dat_in_y1_2, dat_in_y1_1, dat_in_y1_0, dat_in_y0_3, dat_in_y0_2, dat_in_y0_1, dat_in_y0_0 };
  assign dp2reg_lut_hybrid = perf_lut_hybrid_cnt_cur;
  assign dp2reg_lut_le_hit = perf_lut_le_hit_cnt_cur;
  assign dp2reg_lut_lo_hit = perf_lut_lo_hit_cnt_cur;
  assign dp2reg_lut_oflow = perf_lut_oflow_cnt_cur;
  assign dp2reg_lut_uflow = perf_lut_uflow_cnt_cur;
  assign idx2lut_prdy = p1_pipe_ready_bc;
  assign lut_access_type = reg2dp_lut_int_access_type;
  assign lut_addr = reg2dp_lut_int_addr;
  assign lut_data = reg2dp_lut_int_data;
  assign lut_hybrid_cnt = perf_lut_hybrid_cnt_cur;
  assign lut_in_addr0 = p1_pipe_data[288:280];
  assign lut_in_addr0_0 = p1_pipe_data[288:280];
  assign lut_in_addr1 = p1_pipe_data[297:289];
  assign lut_in_addr1_0 = p1_pipe_data[297:289];
  assign lut_in_addr2 = p1_pipe_data[306:298];
  assign lut_in_addr2_0 = p1_pipe_data[306:298];
  assign lut_in_addr3 = p1_pipe_data[315:307];
  assign lut_in_addr3_0 = p1_pipe_data[315:307];
  assign lut_in_fraction0 = p1_pipe_data[34:0];
  assign lut_in_fraction1 = p1_pipe_data[69:35];
  assign lut_in_fraction2 = p1_pipe_data[104:70];
  assign lut_in_fraction3 = p1_pipe_data[139:105];
  assign lut_in_le_hit0 = p1_pipe_data[316];
  assign lut_in_le_hit1 = p1_pipe_data[317];
  assign lut_in_le_hit2 = p1_pipe_data[318];
  assign lut_in_le_hit3 = p1_pipe_data[319];
  assign lut_in_lo_hit0 = p1_pipe_data[320];
  assign lut_in_lo_hit1 = p1_pipe_data[321];
  assign lut_in_lo_hit2 = p1_pipe_data[322];
  assign lut_in_lo_hit3 = p1_pipe_data[323];
  assign lut_in_oflow0 = p1_pipe_data[268];
  assign lut_in_oflow1 = p1_pipe_data[269];
  assign lut_in_oflow2 = p1_pipe_data[270];
  assign lut_in_oflow3 = p1_pipe_data[271];
  assign lut_in_pd = p1_pipe_data;
  assign lut_in_prdy = cmd_fifo_wr_prdy;
  assign lut_in_pvld = p1_pipe_valid;
  assign lut_in_sel0 = p1_pipe_data[276];
  assign lut_in_sel1 = p1_pipe_data[277];
  assign lut_in_sel2 = p1_pipe_data[278];
  assign lut_in_sel3 = p1_pipe_data[279];
  assign lut_in_uflow0 = p1_pipe_data[272];
  assign lut_in_uflow1 = p1_pipe_data[273];
  assign lut_in_uflow2 = p1_pipe_data[274];
  assign lut_in_uflow3 = p1_pipe_data[275];
  assign lut_in_x0 = p1_pipe_data[171:140];
  assign lut_in_x1 = p1_pipe_data[203:172];
  assign lut_in_x2 = p1_pipe_data[235:204];
  assign lut_in_x3 = p1_pipe_data[267:236];
  assign lut_le_hit_cnt = perf_lut_le_hit_cnt_cur;
  assign lut_lo_hit_cnt = perf_lut_lo_hit_cnt_cur;
  assign lut_oflow_cnt = perf_lut_oflow_cnt_cur;
  assign lut_out_pd = { out_flow3, out_flow2, out_flow1, out_flow0, out_bias3, out_bias2, out_bias1, out_bias0, out_offset3, out_offset2, out_offset1, out_offset0, out_shift3, out_shift2, out_shift1, out_shift0, out_scale3, out_scale2, out_scale1, out_scale0, dat_fifo_rd_pd, cmd_fifo_rd_pd[139:0], cmd_fifo_rd_pd[267:140] };
  assign lut_out_prdy = dat_fifo_rd_prdy;
  assign lut_out_pvld = dat_fifo_rd_pvld;
  assign lut_pd = { reg2dp_lut_int_access_type, reg2dp_lut_int_table_id, reg2dp_lut_int_data, reg2dp_lut_int_addr };
  assign lut_table_id = reg2dp_lut_int_table_id;
  assign lut_uflow_cnt = perf_lut_uflow_cnt_cur;
  assign mon_cmd_fifo_rd_pvld = cmd_fifo_rd_pvld;
  assign out_fraction0 = cmd_fifo_rd_pd[34:0];
  assign out_fraction1 = cmd_fifo_rd_pd[69:35];
  assign out_fraction2 = cmd_fifo_rd_pd[104:70];
  assign out_fraction3 = cmd_fifo_rd_pd[139:105];
  assign out_oflow0 = cmd_fifo_rd_pd[268];
  assign out_oflow1 = cmd_fifo_rd_pd[269];
  assign out_oflow2 = cmd_fifo_rd_pd[270];
  assign out_oflow3 = cmd_fifo_rd_pd[271];
  assign out_sel0 = cmd_fifo_rd_pd[276];
  assign out_sel1 = cmd_fifo_rd_pd[277];
  assign out_sel2 = cmd_fifo_rd_pd[278];
  assign out_sel3 = cmd_fifo_rd_pd[279];
  assign out_uflow0 = cmd_fifo_rd_pd[272];
  assign out_uflow1 = cmd_fifo_rd_pd[273];
  assign out_uflow2 = cmd_fifo_rd_pd[274];
  assign out_uflow3 = cmd_fifo_rd_pd[275];
  assign out_x0 = cmd_fifo_rd_pd[171:140];
  assign out_x1 = cmd_fifo_rd_pd[203:172];
  assign out_x2 = cmd_fifo_rd_pd[235:204];
  assign out_x3 = cmd_fifo_rd_pd[267:236];
  assign out_y0_0 = dat_fifo_rd_pd[15:0];
  assign out_y0_1 = dat_fifo_rd_pd[31:16];
  assign out_y0_2 = dat_fifo_rd_pd[47:32];
  assign out_y0_3 = dat_fifo_rd_pd[63:48];
  assign out_y1_0 = dat_fifo_rd_pd[79:64];
  assign out_y1_1 = dat_fifo_rd_pd[95:80];
  assign out_y1_2 = dat_fifo_rd_pd[111:96];
  assign out_y1_3 = dat_fifo_rd_pd[127:112];
  assign p1_assert_clk = nvdla_core_clk;
  assign p1_pipe_rand_data = idx2lut_pd;
  assign p1_pipe_rand_ready = p1_pipe_ready_bc;
  assign p1_pipe_rand_valid = idx2lut_pvld;
  assign p1_pipe_ready = cmd_fifo_wr_prdy;
  assign p2_assert_clk = nvdla_core_clk;
  assign p2_pipe_rand_data = { out_flow3, out_flow2, out_flow1, out_flow0, out_bias3, out_bias2, out_bias1, out_bias0, out_offset3, out_offset2, out_offset1, out_offset0, out_shift3, out_shift2, out_shift1, out_shift0, out_scale3, out_scale2, out_scale1, out_scale0, dat_fifo_rd_pd, cmd_fifo_rd_pd[139:0], cmd_fifo_rd_pd[267:140] };
  assign p2_pipe_rand_ready = dat_fifo_rd_prdy;
  assign p2_pipe_rand_valid = dat_fifo_rd_pvld;
  assign p2_pipe_ready_bc = dat_fifo_rd_prdy;
  assign p2_pipe_skid_data = lut2inp_pd;
  assign p2_pipe_skid_ready = lut2inp_prdy;
  assign p2_pipe_skid_valid = lut2inp_pvld;
  assign p2_skid_ready_flop = p2_pipe_ready;
  assign perf_lut_hybrid_cnt_ext = { 2'b00, perf_lut_hybrid_cnt_cur };
  assign perf_lut_hybrid_sub = 1'b0;
  assign perf_lut_le_hit_cnt_ext = { 2'b00, perf_lut_le_hit_cnt_cur };
  assign perf_lut_le_hit_sub = 1'b0;
  assign perf_lut_lo_hit_cnt_ext = { 2'b00, perf_lut_lo_hit_cnt_cur };
  assign perf_lut_lo_hit_sub = 1'b0;
  assign perf_lut_oflow_cnt_ext = { 2'b00, perf_lut_oflow_cnt_cur };
  assign perf_lut_oflow_sub = 1'b0;
  assign perf_lut_uflow_cnt_ext = { 2'b00, perf_lut_uflow_cnt_cur };
  assign perf_lut_uflow_sub = 1'b0;
  assign pro2lut_pd = { reg2dp_lut_int_access_type, reg2dp_lut_int_table_id, reg2dp_lut_int_data, reg2dp_lut_int_addr };
  assign pro2lut_valid = reg2dp_lut_int_data_wr;
  assign pro_in_addr = reg2dp_lut_int_addr;
  assign pro_in_data = reg2dp_lut_int_data;
  assign pro_in_select_lo = reg2dp_lut_int_table_id;
  assign pro_in_table_id = reg2dp_lut_int_table_id;
  assign pro_in_wr = reg2dp_lut_int_access_type;
  assign rd_lut_en = dat_fifo_wr_pvld;
endmodule
