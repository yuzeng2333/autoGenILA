module \$paramod\SDP_Y_CORE_mgc_io_sync_v1\valid=0 (ld, lz);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:77" *)
  input ld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:78" *)
  output lz;
  assign lz = ld;
endmodule
