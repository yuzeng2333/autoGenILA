module SDP_Y_IDX_leading_sign_32_0(mantissa, rtn);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:144" *)
  wire _000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:158" *)
  wire _001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:158" *)
  wire _002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:159" *)
  wire _003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *)
  wire _004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *)
  wire _005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:165" *)
  wire _006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:168" *)
  wire _007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *)
  wire _008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *)
  wire _009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:170" *)
  wire _010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:171" *)
  wire _011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *)
  wire _012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:136" *)
  wire _029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:143" *)
  wire _030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:149" *)
  wire _031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:157" *)
  wire _032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:132" *)
  wire _033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:133" *)
  wire _034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:134" *)
  wire _035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:138" *)
  wire _036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:139" *)
  wire _037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:140" *)
  wire _038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:145" *)
  wire _039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:146" *)
  wire _040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:147" *)
  wire _041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:151" *)
  wire _042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:152" *)
  wire _043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:153" *)
  wire _044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *)
  wire _045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:161" *)
  wire _053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *)
  wire _054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *)
  wire _055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *)
  wire _056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:165" *)
  wire _057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *)
  wire _058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *)
  wire _059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *)
  wire _060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *)
  wire _063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *)
  wire _064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *)
  wire _065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *)
  wire _085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:161" *)
  wire _086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *)
  wire _087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *)
  wire _088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:167" *)
  wire _089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *)
  wire _090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:171" *)
  wire _091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *)
  wire _092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *)
  wire _093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *)
  wire _094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *)
  wire _096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *)
  wire _097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *)
  wire _098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *)
  wire _100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:125" *)
  wire [4:0] IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:127" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:126" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:128" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:129" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:111" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:103" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:112" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:104" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:113" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:105" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:114" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:106" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:115" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:107" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:110" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:102" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:116" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:108" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:117" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:109" *)
  wire IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:122" *)
  wire c_h_1_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:123" *)
  wire c_h_1_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:124" *)
  wire c_h_1_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:118" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:119" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:120" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:121" *)
  wire c_h_1_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:99" *)
  input [31:0] mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:100" *)
  output [5:0] rtn;
  assign c_h_1_2 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:135" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3 = _029_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:137" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:141" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:142" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _030_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:144" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:144" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:148" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3 = _031_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:150" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1;
  assign c_h_1_12 = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:154" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:155" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:156" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4;
  assign _001_ = _032_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:158" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1;
  assign _002_ = _001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:158" *) c_h_1_12;
  assign _003_ = _002_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:159" *) c_h_1_13;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5 = _003_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:159" *) c_h_1_14;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:161" *) _086_;
  assign _004_ = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *) _087_;
  assign _005_ = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *) _088_;
  assign _006_ = _056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:165" *) c_h_1_14;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl = _004_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:165" *) _057_;
  assign _007_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:168" *) _089_;
  assign _008_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *) _090_;
  assign _009_ = _058_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *) c_h_1_6;
  assign _010_ = _007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:170" *) _059_;
  assign _011_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:171" *) _091_;
  assign _012_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *) _092_;
  assign _013_ = _060_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) c_h_1_13;
  assign _014_ = _011_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) _061_;
  assign _015_ = _062_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) c_h_1_14;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl = _010_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) _063_;
  assign _016_ = _094_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) c_h_1_2;
  assign _017_ = _065_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) _067_;
  assign _018_ = _096_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) c_h_1_5;
  assign _019_ = _069_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _071_;
  assign _020_ = _072_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) c_h_1_6;
  assign _021_ = _017_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _073_;
  assign _022_ = _098_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) c_h_1_9;
  assign _023_ = _075_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) _077_;
  assign _024_ = _100_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) c_h_1_12;
  assign _025_ = _079_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _081_;
  assign _026_ = _082_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) c_h_1_13;
  assign _027_ = _023_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _083_;
  assign _028_ = _084_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) c_h_1_14;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl = _021_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _085_;
  assign _029_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:136" *) mantissa[25:24];
  assign _030_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:143" *) mantissa[17:16];
  assign _031_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:149" *) mantissa[9:8];
  assign _032_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:157" *) mantissa[1:0];
  assign _033_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:132" *) mantissa[29:28];
  assign _034_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:133" *) mantissa[31:30];
  assign _035_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:134" *) mantissa[27:26];
  assign _036_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:138" *) mantissa[21:20];
  assign _037_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:139" *) mantissa[23:22];
  assign _038_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:140" *) mantissa[19:18];
  assign _039_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:145" *) mantissa[13:12];
  assign _040_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:146" *) mantissa[15:14];
  assign _041_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:147" *) mantissa[11:10];
  assign _042_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:151" *) mantissa[5:4];
  assign _043_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:152" *) mantissa[7:6];
  assign _044_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:153" *) mantissa[3:2];
  assign _045_ = mantissa[30:29] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *) 1'b1;
  assign _046_ = mantissa[26:25] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) 1'b1;
  assign _047_ = mantissa[22:21] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) 1'b1;
  assign _048_ = mantissa[18:17] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) 1'b1;
  assign _049_ = mantissa[14:13] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) 1'b1;
  assign _050_ = mantissa[10:9] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) 1'b1;
  assign _051_ = mantissa[6:5] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) 1'b1;
  assign _052_ = mantissa[2:1] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) 1'b1;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:132" *) _033_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:133" *) _034_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:134" *) _035_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:138" *) _036_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:139" *) _037_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:140" *) _038_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:145" *) _039_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:146" *) _040_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:147" *) _041_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:151" *) _042_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_70_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:152" *) _043_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:153" *) _044_;
  assign _053_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:161" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_42_4_sdt_4;
  assign _054_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_18_3_sdt_3;
  assign _055_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *) IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_62_3_sdt_3;
  assign _056_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *) _005_;
  assign _057_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:165" *) _006_;
  assign _058_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *) _008_;
  assign _059_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *) _009_;
  assign _060_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *) _012_;
  assign _061_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) _013_;
  assign _062_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) _014_;
  assign _063_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:173" *) _015_;
  assign _064_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *) _045_;
  assign _065_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *) _093_;
  assign _066_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) _046_;
  assign _067_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) _016_;
  assign _068_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) _047_;
  assign _069_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) _095_;
  assign _070_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) _048_;
  assign _071_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _018_;
  assign _072_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _019_;
  assign _073_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _020_;
  assign _074_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _049_;
  assign _075_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _097_;
  assign _076_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) _050_;
  assign _077_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) _022_;
  assign _078_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) _051_;
  assign _079_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) _099_;
  assign _080_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) _052_;
  assign _081_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _024_;
  assign _082_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _025_;
  assign _083_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _026_;
  assign _084_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _027_;
  assign _085_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:180" *) _028_;
  assign _086_ = c_h_1_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:161" *) _053_;
  assign _087_ = c_h_1_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:163" *) _054_;
  assign _088_ = c_h_1_12 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:164" *) _055_;
  assign _089_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:167" *) _033_;
  assign _090_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:169" *) _036_;
  assign _091_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_58_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:171" *) _039_;
  assign _092_ = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_78_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:172" *) _042_;
  assign _093_ = mantissa[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:174" *) _064_;
  assign _094_ = mantissa[27] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:175" *) _066_;
  assign _095_ = mantissa[23] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) _068_;
  assign _096_ = mantissa[19] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:176" *) _070_;
  assign _097_ = mantissa[15] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:177" *) _074_;
  assign _098_ = mantissa[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:178" *) _076_;
  assign _099_ = mantissa[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) _078_;
  assign _100_ = mantissa[3] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:179" *) _080_;
  assign IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl = IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:194|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:193" *) 5'b00000 : { c_h_1_14, IntLeadZero_32U_leading_sign_32_0_rtn_and_119_nl, IntLeadZero_32U_leading_sign_32_0_rtn_and_117_nl, IntLeadZero_32U_leading_sign_32_0_rtn_and_124_nl, IntLeadZero_32U_leading_sign_32_0_rtn_and_127_nl };
  assign rtn = { IntLeadZero_32U_leading_sign_32_0_rtn_wrs_c_92_5_sdt_5, IntLeadZero_32U_leading_sign_32_0_rtn_IntLeadZero_32U_leading_sign_32_0_rtn_and_nl };
endmodule
