module CDP_OCVT_chn_data_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:273" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:274" *)
  output outsig;
  assign outsig = in_0;
endmodule
