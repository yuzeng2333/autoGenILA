module aes_top(clk, rst, wr, addr, data_in, data_out, ack, stb, xram_addr, xram_data_out, xram_data_in, xram_ack, xram_stb, xram_wr, aes_state, aes_addr, aes_len, aes_ctr, aes_key0, aes_step);
  logic [1:0] _000_;
  logic [4:0] _001_;
  logic [15:0] _002_;
  logic [3:0] _003_;
  logic [127:0] _004_;
  logic [127:0] _005_;
  logic [15:0] _006_;
  logic [127:0] _007_;
  logic [15:0] _008_;
  logic [15:0] _009_;
  logic [3:0] _010_;
  logic [15:0] _011_;
  logic [127:0] _012_;
  logic [4:0] _013_;
  logic [31:0] _014_;
  logic _015_;
  logic _016_;
  logic _017_;
  logic _018_;
  logic _019_;
  logic _020_;
  logic _021_;
  logic _022_;
  logic _023_;
  logic _024_;
  logic _025_;
  logic _026_;
  logic _027_;
  logic _028_;
  logic _029_;
  logic _030_;
  logic _031_;
  logic _032_;
  logic _033_;
  logic _034_;
  logic _035_;
  logic _036_;
  logic _037_;
  logic _038_;
  logic _039_;
  logic _040_;
  logic _041_;
  logic _042_;
  logic _043_;
  logic _044_;
  logic _045_;
  logic _046_;
  logic _047_;
  logic _048_;
  logic _049_;
  logic _050_;
  logic _051_;
  logic _052_;
  logic _053_;
  logic [127:0] _054_;
  logic _055_;
  logic _056_;
  logic _057_;
  logic _058_;
  logic _059_;
  logic _060_;
  logic _061_;
  logic _062_;
  logic _063_;
  logic _064_;
  logic _065_;
  logic _066_;
  logic _067_;
  logic _068_;
  logic _069_;
  logic _070_;
  logic _071_;
  logic [7:0] _072_;
  logic [7:0] _073_;
  logic [7:0] _074_;
  logic [7:0] _075_;
  logic [7:0] _076_;
  logic [7:0] _077_;
  logic [7:0] _078_;
  logic [7:0] _079_;
  logic [7:0] _080_;
  logic [7:0] _081_;
  logic [7:0] _082_;
  logic [7:0] _083_;
  logic [7:0] _084_;
  logic [7:0] _085_;
  logic [127:0] _086_;
  logic _087_;
  logic [7:0] _088_;
  logic [7:0] _089_;
  logic [7:0] _090_;
  logic [7:0] _091_;
  logic [7:0] _092_;
  logic [7:0] _093_;
  logic [7:0] _094_;
  logic [7:0] _095_;
  logic [7:0] _096_;
  logic [7:0] _097_;
  logic [7:0] _098_;
  logic [7:0] _099_;
  logic [7:0] _100_;
  logic [7:0] _101_;
  logic [15:0] _102_;
  logic _103_;
  logic _104_;
  logic [15:0] _105_;
  logic _106_;
  logic [7:0] _107_;
  logic [7:0] _108_;
  logic [7:0] _109_;
  logic [7:0] _110_;
  logic [31:0] _111_;
  logic [31:0] _112_;
  logic [1:0] _113_;
  logic [1:0] _114_;
  logic [1:0] _115_;
  logic [1:0] _116_;
  logic [127:0] _117_;
  logic [4:0] _118_;
  logic [7:0] _119_;
  logic [7:0] _120_;
  logic [7:0] _121_;
  logic [7:0] _122_;
  logic [7:0] _123_;
  logic [7:0] _124_;
  logic [7:0] _125_;
  logic [7:0] _126_;
  logic [7:0] _127_;
  logic [7:0] _128_;
  logic [7:0] _129_;
  logic [7:0] _130_;
  logic [7:0] _131_;
  logic [7:0] _132_;
  output ack;
  input [15:0] addr;
  output [15:0] aes_addr;
  logic [7:0] aes_addr_dataout;
  output [127:0] aes_ctr;
  logic [7:0] aes_ctr_dataout;
  logic [127:0] aes_curr_key;
  output [127:0] aes_key0;
  logic [7:0] aes_key0_dataout;
  output [15:0] aes_len;
  logic [7:0] aes_len_dataout;
  logic [127:0] aes_out;
  logic [127:0] aes_reg_ctr;
  logic [3:0] \aes_reg_ctr_i.addr ;
  logic \aes_reg_ctr_i.clk ;
  logic [7:0] \aes_reg_ctr_i.data_in ;
  logic [7:0] \aes_reg_ctr_i.data_out ;
  logic [7:0] \aes_reg_ctr_i.data_out_mux ;
  logic \aes_reg_ctr_i.en ;
  logic [7:0] \aes_reg_ctr_i.reg0_next ;
  logic [7:0] \aes_reg_ctr_i.reg10_next ;
  logic [7:0] \aes_reg_ctr_i.reg11_next ;
  logic [7:0] \aes_reg_ctr_i.reg12_next ;
  logic [7:0] \aes_reg_ctr_i.reg13_next ;
  logic [7:0] \aes_reg_ctr_i.reg14_next ;
  logic [7:0] \aes_reg_ctr_i.reg15_next ;
  logic [7:0] \aes_reg_ctr_i.reg1_next ;
  logic [7:0] \aes_reg_ctr_i.reg2_next ;
  logic [7:0] \aes_reg_ctr_i.reg3_next ;
  logic [7:0] \aes_reg_ctr_i.reg4_next ;
  logic [7:0] \aes_reg_ctr_i.reg5_next ;
  logic [7:0] \aes_reg_ctr_i.reg6_next ;
  logic [7:0] \aes_reg_ctr_i.reg7_next ;
  logic [7:0] \aes_reg_ctr_i.reg8_next ;
  logic [7:0] \aes_reg_ctr_i.reg9_next ;
  logic [127:0] \aes_reg_ctr_i.reg_out ;
  logic \aes_reg_ctr_i.rst ;
  logic \aes_reg_ctr_i.wr ;
  logic \aes_reg_ctr_i.wr0 ;
  logic \aes_reg_ctr_i.wr1 ;
  logic \aes_reg_ctr_i.wr10 ;
  logic \aes_reg_ctr_i.wr11 ;
  logic \aes_reg_ctr_i.wr12 ;
  logic \aes_reg_ctr_i.wr13 ;
  logic \aes_reg_ctr_i.wr14 ;
  logic \aes_reg_ctr_i.wr15 ;
  logic \aes_reg_ctr_i.wr2 ;
  logic \aes_reg_ctr_i.wr3 ;
  logic \aes_reg_ctr_i.wr4 ;
  logic \aes_reg_ctr_i.wr5 ;
  logic \aes_reg_ctr_i.wr6 ;
  logic \aes_reg_ctr_i.wr7 ;
  logic \aes_reg_ctr_i.wr8 ;
  logic \aes_reg_ctr_i.wr9 ;
  logic [127:0] aes_reg_key0;
  logic [3:0] \aes_reg_key0_i.addr ;
  logic \aes_reg_key0_i.clk ;
  logic [7:0] \aes_reg_key0_i.data_in ;
  logic [7:0] \aes_reg_key0_i.data_out ;
  logic [7:0] \aes_reg_key0_i.data_out_mux ;
  logic \aes_reg_key0_i.en ;
  logic [7:0] \aes_reg_key0_i.reg0_next ;
  logic [7:0] \aes_reg_key0_i.reg10_next ;
  logic [7:0] \aes_reg_key0_i.reg11_next ;
  logic [7:0] \aes_reg_key0_i.reg12_next ;
  logic [7:0] \aes_reg_key0_i.reg13_next ;
  logic [7:0] \aes_reg_key0_i.reg14_next ;
  logic [7:0] \aes_reg_key0_i.reg15_next ;
  logic [7:0] \aes_reg_key0_i.reg1_next ;
  logic [7:0] \aes_reg_key0_i.reg2_next ;
  logic [7:0] \aes_reg_key0_i.reg3_next ;
  logic [7:0] \aes_reg_key0_i.reg4_next ;
  logic [7:0] \aes_reg_key0_i.reg5_next ;
  logic [7:0] \aes_reg_key0_i.reg6_next ;
  logic [7:0] \aes_reg_key0_i.reg7_next ;
  logic [7:0] \aes_reg_key0_i.reg8_next ;
  logic [7:0] \aes_reg_key0_i.reg9_next ;
  logic [127:0] \aes_reg_key0_i.reg_out ;
  logic \aes_reg_key0_i.rst ;
  logic \aes_reg_key0_i.wr ;
  logic \aes_reg_key0_i.wr0 ;
  logic \aes_reg_key0_i.wr1 ;
  logic \aes_reg_key0_i.wr10 ;
  logic \aes_reg_key0_i.wr11 ;
  logic \aes_reg_key0_i.wr12 ;
  logic \aes_reg_key0_i.wr13 ;
  logic \aes_reg_key0_i.wr14 ;
  logic \aes_reg_key0_i.wr15 ;
  logic \aes_reg_key0_i.wr2 ;
  logic \aes_reg_key0_i.wr3 ;
  logic \aes_reg_key0_i.wr4 ;
  logic \aes_reg_key0_i.wr5 ;
  logic \aes_reg_key0_i.wr6 ;
  logic \aes_reg_key0_i.wr7 ;
  logic \aes_reg_key0_i.wr8 ;
  logic \aes_reg_key0_i.wr9 ;
  logic [15:0] aes_reg_opaddr;
  logic \aes_reg_opaddr_i.addr ;
  logic \aes_reg_opaddr_i.clk ;
  logic [7:0] \aes_reg_opaddr_i.data_in ;
  logic [7:0] \aes_reg_opaddr_i.data_out ;
  logic [7:0] \aes_reg_opaddr_i.data_out_mux ;
  logic \aes_reg_opaddr_i.en ;
  logic [7:0] \aes_reg_opaddr_i.reg0_next ;
  logic [7:0] \aes_reg_opaddr_i.reg1_next ;
  logic [15:0] \aes_reg_opaddr_i.reg_out ;
  logic \aes_reg_opaddr_i.rst ;
  logic \aes_reg_opaddr_i.wr ;
  logic \aes_reg_opaddr_i.wr0 ;
  logic \aes_reg_opaddr_i.wr1 ;
  logic [15:0] aes_reg_oplen;
  logic \aes_reg_oplen_i.addr ;
  logic \aes_reg_oplen_i.clk ;
  logic [7:0] \aes_reg_oplen_i.data_in ;
  logic [7:0] \aes_reg_oplen_i.data_out ;
  logic [7:0] \aes_reg_oplen_i.data_out_mux ;
  logic \aes_reg_oplen_i.en ;
  logic [7:0] \aes_reg_oplen_i.reg0_next ;
  logic [7:0] \aes_reg_oplen_i.reg1_next ;
  logic [15:0] \aes_reg_oplen_i.reg_out ;
  logic \aes_reg_oplen_i.rst ;
  logic \aes_reg_oplen_i.wr ;
  logic \aes_reg_oplen_i.wr0 ;
  logic \aes_reg_oplen_i.wr1 ;
  logic [1:0] aes_reg_state;
  logic [1:0] aes_reg_state_next;
  logic aes_reg_state_next_idle;
  logic aes_reg_state_next_operate;
  logic [1:0] aes_reg_state_next_read_data;
  logic [1:0] aes_reg_state_next_write_data;
  output [1:0] aes_state;
  logic aes_state_idle;
  logic aes_state_operate;
  logic aes_state_read_data;
  logic aes_state_write_data;
  output aes_step;
  logic [4:0] aes_time_counter;
  logic [4:0] aes_time_counter_next;
  logic aes_time_enough;
  logic [15:0] block_counter;
  logic [15:0] block_counter_next;
  logic [3:0] byte_counter;
  logic [3:0] byte_counter_next;
  input clk;
  input [7:0] data_in;
  output [7:0] data_out;
  logic [127:0] encrypted_data;
  logic [127:0] encrypted_data_buf;
  logic [127:0] encrypted_data_buf_next;
  logic in_addr_range;
  logic incr_byte_counter;
  logic last_byte_acked;
  logic [127:0] mem_data_buf;
  logic [127:0] mem_data_buf_next;
  logic more_blocks;
  logic [15:0] operated_bytes_count;
  logic [15:0] operated_bytes_count_next;
  logic reset_byte_counter;
  input rst;
  logic sel_reg_addr;
  logic sel_reg_ctr;
  logic sel_reg_key0;
  logic sel_reg_len;
  logic sel_reg_start;
  logic sel_reg_state;
  logic start_op;
  input stb;
  logic [127:0] uaes_ctr;
  logic [127:0] uaes_ctr_nxt;
  input wr;
  logic wren;
  input xram_ack;
  output [15:0] xram_addr;
  input [7:0] xram_data_in;
  output [7:0] xram_data_out;
  output xram_stb;
  output xram_wr;
  assign _008_ = operated_bytes_count + 5'b10000;
  assign _009_ = block_counter + 5'b10000;
  assign _010_ = byte_counter + 1'b1;
  assign _011_ = \aes_reg_opaddr_i.reg_out + block_counter;
  assign xram_addr = _011_ + byte_counter;
  assign _012_ = uaes_ctr + 5'b10000;
  assign _013_ = aes_time_counter + 1'b1;
  assign sel_reg_start = addr == 16'b1111111100000000;
  assign sel_reg_state = addr == 16'b1111111100000001;
  assign \aes_reg_opaddr_i.en = addr[15:1] == 15'b111111110000001;
  assign \aes_reg_oplen_i.en = addr[15:1] == 15'b111111110000010;
  assign \aes_reg_ctr_i.en = addr[15:4] == 12'b111111110010;
  assign \aes_reg_key0_i.en = addr[15:4] == 12'b111111110001;
  assign aes_state_idle = ! aes_reg_state;
  assign aes_state_read_data = aes_reg_state == 1'b1;
  assign aes_state_operate = aes_reg_state == 2'b10;
  assign aes_state_write_data = aes_reg_state == 2'b11;
  assign _015_ = byte_counter == 4'b1111;
  assign _016_ = ! byte_counter;
  assign _017_ = byte_counter == 1'b1;
  assign _018_ = byte_counter == 2'b10;
  assign _019_ = byte_counter == 2'b11;
  assign _020_ = byte_counter == 3'b100;
  assign _021_ = byte_counter == 3'b101;
  assign _022_ = byte_counter == 3'b110;
  assign _023_ = byte_counter == 3'b111;
  assign _024_ = byte_counter == 4'b1000;
  assign _025_ = byte_counter == 4'b1001;
  assign _026_ = byte_counter == 4'b1010;
  assign _027_ = byte_counter == 4'b1011;
  assign _028_ = byte_counter == 4'b1100;
  assign _029_ = byte_counter == 4'b1101;
  assign _030_ = byte_counter == 4'b1110;
  assign _031_ = addr >= 16'b1111111100000000;
  assign aes_time_enough = aes_time_counter >= 5'b10100;
  assign in_addr_range = _031_ && _051_;
  assign ack = stb && in_addr_range;
  assign wren = wr && aes_state_idle;
  assign _032_ = sel_reg_start && data_in[0];
  assign reset_byte_counter = _032_ && wren;
  assign \aes_reg_opaddr_i.wr = \aes_reg_opaddr_i.en && wren;
  assign \aes_reg_oplen_i.wr = \aes_reg_oplen_i.en && wren;
  assign \aes_reg_ctr_i.wr = \aes_reg_ctr_i.en && wren;
  assign \aes_reg_key0_i.wr = \aes_reg_key0_i.en && wren;
  assign _033_ = last_byte_acked && aes_state_write_data;
  assign last_byte_acked = _015_ && xram_ack;
  assign more_blocks = _033_ && _052_;
  assign _034_ = last_byte_acked && more_blocks;
  assign _035_ = xram_ack && _016_;
  assign _036_ = xram_ack && _017_;
  assign _037_ = xram_ack && _018_;
  assign _038_ = xram_ack && _019_;
  assign _039_ = xram_ack && _020_;
  assign _040_ = xram_ack && _021_;
  assign _041_ = xram_ack && _022_;
  assign _042_ = xram_ack && _023_;
  assign _043_ = xram_ack && _024_;
  assign _044_ = xram_ack && _025_;
  assign _045_ = xram_ack && _026_;
  assign _046_ = xram_ack && _027_;
  assign _047_ = xram_ack && _028_;
  assign _048_ = xram_ack && _029_;
  assign _049_ = xram_ack && _030_;
  assign xram_stb = aes_state_read_data || aes_state_write_data;
  assign _050_ = more_blocks || reset_byte_counter;
  assign _051_ = addr < 16'b1111111100110000;
  assign _052_ = operated_bytes_count_next < \aes_reg_oplen_i.reg_out ;
  assign _053_ = aes_time_counter < 5'b11111;
  assign aes_step = aes_reg_state != aes_reg_state_next;
  always @(posedge clk)
      aes_reg_state <= _000_;
  always @(posedge clk)
      operated_bytes_count <= _006_;
  always @(posedge clk)
      block_counter <= _002_;
  always @(posedge clk)
      byte_counter <= _003_;
  always @(posedge clk)
      mem_data_buf <= _005_;
  always @(posedge clk)
      encrypted_data_buf <= _004_;
  always @(posedge clk)
      aes_time_counter <= _001_;
  always @(posedge clk)
      uaes_ctr <= _007_;
  assign _004_ = rst ? encrypted_data_buf : encrypted_data_buf_next;
  assign _005_ = rst ? mem_data_buf : mem_data_buf_next;
  assign _003_ = rst ? 4'b0000 : byte_counter_next;
  assign _002_ = rst ? 16'b0000000000000000 : block_counter_next;
  assign _006_ = rst ? 16'b0000000000000000 : operated_bytes_count_next;
  assign _000_ = rst ? 2'b00 : aes_reg_state_next;
  assign _001_ = rst ? 5'b00000 : aes_time_counter_next;
  assign _007_ = rst ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : uaes_ctr_nxt;
  assign _055_ = ! addr[3:0];
  assign _056_ = addr[3:0] == 1'b1;
  assign _057_ = addr[3:0] == 2'b10;
  assign _058_ = addr[3:0] == 2'b11;
  assign _059_ = addr[3:0] == 3'b100;
  assign _060_ = addr[3:0] == 3'b101;
  assign _061_ = addr[3:0] == 3'b110;
  assign _062_ = addr[3:0] == 3'b111;
  assign _063_ = addr[3:0] == 4'b1000;
  assign _064_ = addr[3:0] == 4'b1001;
  assign _065_ = addr[3:0] == 4'b1010;
  assign _066_ = addr[3:0] == 4'b1011;
  assign _067_ = addr[3:0] == 4'b1100;
  assign _068_ = addr[3:0] == 4'b1101;
  assign _069_ = addr[3:0] == 4'b1110;
  assign _070_ = addr[3:0] == 4'b1111;
  assign _071_ = \aes_reg_ctr_i.en && \aes_reg_ctr_i.wr ;
  assign \aes_reg_ctr_i.wr0 = _071_ && _055_;
  assign \aes_reg_ctr_i.wr1 = _071_ && _056_;
  assign \aes_reg_ctr_i.wr2 = _071_ && _057_;
  assign \aes_reg_ctr_i.wr3 = _071_ && _058_;
  assign \aes_reg_ctr_i.wr4 = _071_ && _059_;
  assign \aes_reg_ctr_i.wr5 = _071_ && _060_;
  assign \aes_reg_ctr_i.wr6 = _071_ && _061_;
  assign \aes_reg_ctr_i.wr7 = _071_ && _062_;
  assign \aes_reg_ctr_i.wr8 = _071_ && _063_;
  assign \aes_reg_ctr_i.wr9 = _071_ && _064_;
  assign \aes_reg_ctr_i.wr10 = _071_ && _065_;
  assign \aes_reg_ctr_i.wr11 = _071_ && _066_;
  assign \aes_reg_ctr_i.wr12 = _071_ && _067_;
  assign \aes_reg_ctr_i.wr13 = _071_ && _068_;
  assign \aes_reg_ctr_i.wr14 = _071_ && _069_;
  assign \aes_reg_ctr_i.wr15 = _071_ && _070_;
  always @(posedge clk)
      \aes_reg_ctr_i.reg_out <= _054_;
  assign _054_[127:120] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg15_next ;
  assign _054_[119:112] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg14_next ;
  assign _054_[111:104] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg13_next ;
  assign _054_[103:96] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg12_next ;
  assign _054_[95:88] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg11_next ;
  assign _054_[87:80] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg10_next ;
  assign _054_[79:72] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg9_next ;
  assign _054_[71:64] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg8_next ;
  assign _054_[63:56] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg7_next ;
  assign _054_[55:48] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg6_next ;
  assign _054_[47:40] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg5_next ;
  assign _054_[39:32] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg4_next ;
  assign _054_[31:24] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg3_next ;
  assign _054_[23:16] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg2_next ;
  assign _054_[15:8] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg1_next ;
  assign _054_[7:0] = rst ? 8'b00000000 : \aes_reg_ctr_i.reg0_next ;
  assign \aes_reg_ctr_i.reg0_next = \aes_reg_ctr_i.wr0 ? data_in : \aes_reg_ctr_i.reg_out [7:0];
  assign \aes_reg_ctr_i.reg1_next = \aes_reg_ctr_i.wr1 ? data_in : \aes_reg_ctr_i.reg_out [15:8];
  assign \aes_reg_ctr_i.reg2_next = \aes_reg_ctr_i.wr2 ? data_in : \aes_reg_ctr_i.reg_out [23:16];
  assign \aes_reg_ctr_i.reg3_next = \aes_reg_ctr_i.wr3 ? data_in : \aes_reg_ctr_i.reg_out [31:24];
  assign \aes_reg_ctr_i.reg4_next = \aes_reg_ctr_i.wr4 ? data_in : \aes_reg_ctr_i.reg_out [39:32];
  assign \aes_reg_ctr_i.reg5_next = \aes_reg_ctr_i.wr5 ? data_in : \aes_reg_ctr_i.reg_out [47:40];
  assign \aes_reg_ctr_i.reg6_next = \aes_reg_ctr_i.wr6 ? data_in : \aes_reg_ctr_i.reg_out [55:48];
  assign \aes_reg_ctr_i.reg7_next = \aes_reg_ctr_i.wr7 ? data_in : \aes_reg_ctr_i.reg_out [63:56];
  assign \aes_reg_ctr_i.reg8_next = \aes_reg_ctr_i.wr8 ? data_in : \aes_reg_ctr_i.reg_out [71:64];
  assign \aes_reg_ctr_i.reg9_next = \aes_reg_ctr_i.wr9 ? data_in : \aes_reg_ctr_i.reg_out [79:72];
  assign \aes_reg_ctr_i.reg10_next = \aes_reg_ctr_i.wr10 ? data_in : \aes_reg_ctr_i.reg_out [87:80];
  assign \aes_reg_ctr_i.reg11_next = \aes_reg_ctr_i.wr11 ? data_in : \aes_reg_ctr_i.reg_out [95:88];
  assign \aes_reg_ctr_i.reg12_next = \aes_reg_ctr_i.wr12 ? data_in : \aes_reg_ctr_i.reg_out [103:96];
  assign \aes_reg_ctr_i.reg13_next = \aes_reg_ctr_i.wr13 ? data_in : \aes_reg_ctr_i.reg_out [111:104];
  assign \aes_reg_ctr_i.reg14_next = \aes_reg_ctr_i.wr14 ? data_in : \aes_reg_ctr_i.reg_out [119:112];
  assign \aes_reg_ctr_i.reg15_next = \aes_reg_ctr_i.wr15 ? data_in : \aes_reg_ctr_i.reg_out [127:120];
  assign _072_ = _069_ ? \aes_reg_ctr_i.reg_out [119:112] : \aes_reg_ctr_i.reg_out [127:120];
  assign _073_ = _068_ ? \aes_reg_ctr_i.reg_out [111:104] : _072_;
  assign _074_ = _067_ ? \aes_reg_ctr_i.reg_out [103:96] : _073_;
  assign _075_ = _066_ ? \aes_reg_ctr_i.reg_out [95:88] : _074_;
  assign _076_ = _065_ ? \aes_reg_ctr_i.reg_out [87:80] : _075_;
  assign _077_ = _064_ ? \aes_reg_ctr_i.reg_out [79:72] : _076_;
  assign _078_ = _063_ ? \aes_reg_ctr_i.reg_out [71:64] : _077_;
  assign _079_ = _062_ ? \aes_reg_ctr_i.reg_out [63:56] : _078_;
  assign _080_ = _061_ ? \aes_reg_ctr_i.reg_out [55:48] : _079_;
  assign _081_ = _060_ ? \aes_reg_ctr_i.reg_out [47:40] : _080_;
  assign _082_ = _059_ ? \aes_reg_ctr_i.reg_out [39:32] : _081_;
  assign _083_ = _058_ ? \aes_reg_ctr_i.reg_out [31:24] : _082_;
  assign _084_ = _057_ ? \aes_reg_ctr_i.reg_out [23:16] : _083_;
  assign _085_ = _056_ ? \aes_reg_ctr_i.reg_out [15:8] : _084_;
  assign aes_ctr_dataout = _055_ ? \aes_reg_ctr_i.reg_out [7:0] : _085_;
  assign _087_ = \aes_reg_key0_i.en && \aes_reg_key0_i.wr ;
  assign \aes_reg_key0_i.wr0 = _087_ && _055_;
  assign \aes_reg_key0_i.wr1 = _087_ && _056_;
  assign \aes_reg_key0_i.wr2 = _087_ && _057_;
  assign \aes_reg_key0_i.wr3 = _087_ && _058_;
  assign \aes_reg_key0_i.wr4 = _087_ && _059_;
  assign \aes_reg_key0_i.wr5 = _087_ && _060_;
  assign \aes_reg_key0_i.wr6 = _087_ && _061_;
  assign \aes_reg_key0_i.wr7 = _087_ && _062_;
  assign \aes_reg_key0_i.wr8 = _087_ && _063_;
  assign \aes_reg_key0_i.wr9 = _087_ && _064_;
  assign \aes_reg_key0_i.wr10 = _087_ && _065_;
  assign \aes_reg_key0_i.wr11 = _087_ && _066_;
  assign \aes_reg_key0_i.wr12 = _087_ && _067_;
  assign \aes_reg_key0_i.wr13 = _087_ && _068_;
  assign \aes_reg_key0_i.wr14 = _087_ && _069_;
  assign \aes_reg_key0_i.wr15 = _087_ && _070_;
  always @(posedge clk)
      \aes_reg_key0_i.reg_out <= _086_;
  assign _086_[127:120] = rst ? 8'b00000000 : \aes_reg_key0_i.reg15_next ;
  assign _086_[119:112] = rst ? 8'b00000000 : \aes_reg_key0_i.reg14_next ;
  assign _086_[111:104] = rst ? 8'b00000000 : \aes_reg_key0_i.reg13_next ;
  assign _086_[103:96] = rst ? 8'b00000000 : \aes_reg_key0_i.reg12_next ;
  assign _086_[95:88] = rst ? 8'b00000000 : \aes_reg_key0_i.reg11_next ;
  assign _086_[87:80] = rst ? 8'b00000000 : \aes_reg_key0_i.reg10_next ;
  assign _086_[79:72] = rst ? 8'b00000000 : \aes_reg_key0_i.reg9_next ;
  assign _086_[71:64] = rst ? 8'b00000000 : \aes_reg_key0_i.reg8_next ;
  assign _086_[63:56] = rst ? 8'b00000000 : \aes_reg_key0_i.reg7_next ;
  assign _086_[55:48] = rst ? 8'b00000000 : \aes_reg_key0_i.reg6_next ;
  assign _086_[47:40] = rst ? 8'b00000000 : \aes_reg_key0_i.reg5_next ;
  assign _086_[39:32] = rst ? 8'b00000000 : \aes_reg_key0_i.reg4_next ;
  assign _086_[31:24] = rst ? 8'b00000000 : \aes_reg_key0_i.reg3_next ;
  assign _086_[23:16] = rst ? 8'b00000000 : \aes_reg_key0_i.reg2_next ;
  assign _086_[15:8] = rst ? 8'b00000000 : \aes_reg_key0_i.reg1_next ;
  assign _086_[7:0] = rst ? 8'b00000000 : \aes_reg_key0_i.reg0_next ;
  assign \aes_reg_key0_i.reg0_next = \aes_reg_key0_i.wr0 ? data_in : \aes_reg_key0_i.reg_out [7:0];
  assign \aes_reg_key0_i.reg1_next = \aes_reg_key0_i.wr1 ? data_in : \aes_reg_key0_i.reg_out [15:8];
  assign \aes_reg_key0_i.reg2_next = \aes_reg_key0_i.wr2 ? data_in : \aes_reg_key0_i.reg_out [23:16];
  assign \aes_reg_key0_i.reg3_next = \aes_reg_key0_i.wr3 ? data_in : \aes_reg_key0_i.reg_out [31:24];
  assign \aes_reg_key0_i.reg4_next = \aes_reg_key0_i.wr4 ? data_in : \aes_reg_key0_i.reg_out [39:32];
  assign \aes_reg_key0_i.reg5_next = \aes_reg_key0_i.wr5 ? data_in : \aes_reg_key0_i.reg_out [47:40];
  assign \aes_reg_key0_i.reg6_next = \aes_reg_key0_i.wr6 ? data_in : \aes_reg_key0_i.reg_out [55:48];
  assign \aes_reg_key0_i.reg7_next = \aes_reg_key0_i.wr7 ? data_in : \aes_reg_key0_i.reg_out [63:56];
  assign \aes_reg_key0_i.reg8_next = \aes_reg_key0_i.wr8 ? data_in : \aes_reg_key0_i.reg_out [71:64];
  assign \aes_reg_key0_i.reg9_next = \aes_reg_key0_i.wr9 ? data_in : \aes_reg_key0_i.reg_out [79:72];
  assign \aes_reg_key0_i.reg10_next = \aes_reg_key0_i.wr10 ? data_in : \aes_reg_key0_i.reg_out [87:80];
  assign \aes_reg_key0_i.reg11_next = \aes_reg_key0_i.wr11 ? data_in : \aes_reg_key0_i.reg_out [95:88];
  assign \aes_reg_key0_i.reg12_next = \aes_reg_key0_i.wr12 ? data_in : \aes_reg_key0_i.reg_out [103:96];
  assign \aes_reg_key0_i.reg13_next = \aes_reg_key0_i.wr13 ? data_in : \aes_reg_key0_i.reg_out [111:104];
  assign \aes_reg_key0_i.reg14_next = \aes_reg_key0_i.wr14 ? data_in : \aes_reg_key0_i.reg_out [119:112];
  assign \aes_reg_key0_i.reg15_next = \aes_reg_key0_i.wr15 ? data_in : \aes_reg_key0_i.reg_out [127:120];
  assign _088_ = _069_ ? \aes_reg_key0_i.reg_out [119:112] : \aes_reg_key0_i.reg_out [127:120];
  assign _089_ = _068_ ? \aes_reg_key0_i.reg_out [111:104] : _088_;
  assign _090_ = _067_ ? \aes_reg_key0_i.reg_out [103:96] : _089_;
  assign _091_ = _066_ ? \aes_reg_key0_i.reg_out [95:88] : _090_;
  assign _092_ = _065_ ? \aes_reg_key0_i.reg_out [87:80] : _091_;
  assign _093_ = _064_ ? \aes_reg_key0_i.reg_out [79:72] : _092_;
  assign _094_ = _063_ ? \aes_reg_key0_i.reg_out [71:64] : _093_;
  assign _095_ = _062_ ? \aes_reg_key0_i.reg_out [63:56] : _094_;
  assign _096_ = _061_ ? \aes_reg_key0_i.reg_out [55:48] : _095_;
  assign _097_ = _060_ ? \aes_reg_key0_i.reg_out [47:40] : _096_;
  assign _098_ = _059_ ? \aes_reg_key0_i.reg_out [39:32] : _097_;
  assign _099_ = _058_ ? \aes_reg_key0_i.reg_out [31:24] : _098_;
  assign _100_ = _057_ ? \aes_reg_key0_i.reg_out [23:16] : _099_;
  assign _101_ = _056_ ? \aes_reg_key0_i.reg_out [15:8] : _100_;
  assign aes_key0_dataout = _055_ ? \aes_reg_key0_i.reg_out [7:0] : _101_;
  assign _103_ = ~ addr[0];
  assign _104_ = \aes_reg_opaddr_i.en && \aes_reg_opaddr_i.wr ;
  assign \aes_reg_opaddr_i.wr0 = _104_ && _103_;
  assign \aes_reg_opaddr_i.wr1 = _104_ && addr[0];
  always @(posedge clk)
      \aes_reg_opaddr_i.reg_out <= _102_;
  assign _102_[15:8] = rst ? 8'b00000000 : \aes_reg_opaddr_i.reg1_next ;
  assign _102_[7:0] = rst ? 8'b00000000 : \aes_reg_opaddr_i.reg0_next ;
  assign \aes_reg_opaddr_i.reg0_next = \aes_reg_opaddr_i.wr0 ? data_in : \aes_reg_opaddr_i.reg_out [7:0];
  assign \aes_reg_opaddr_i.reg1_next = \aes_reg_opaddr_i.wr1 ? data_in : \aes_reg_opaddr_i.reg_out [15:8];
  assign aes_addr_dataout = addr[0] ? \aes_reg_opaddr_i.reg_out [15:8] : \aes_reg_opaddr_i.reg_out [7:0];
  assign _106_ = \aes_reg_oplen_i.en && \aes_reg_oplen_i.wr ;
  assign \aes_reg_oplen_i.wr0 = _106_ && _103_;
  assign \aes_reg_oplen_i.wr1 = _106_ && addr[0];
  always @(posedge clk)
      \aes_reg_oplen_i.reg_out <= _105_;
  assign _105_[15:8] = rst ? 8'b00000000 : \aes_reg_oplen_i.reg1_next ;
  assign _105_[7:0] = rst ? 8'b00000000 : \aes_reg_oplen_i.reg0_next ;
  assign \aes_reg_oplen_i.reg0_next = \aes_reg_oplen_i.wr0 ? data_in : \aes_reg_oplen_i.reg_out [7:0];
  assign \aes_reg_oplen_i.reg1_next = \aes_reg_oplen_i.wr1 ? data_in : \aes_reg_oplen_i.reg_out [15:8];
  assign aes_len_dataout = addr[0] ? \aes_reg_oplen_i.reg_out [15:8] : \aes_reg_oplen_i.reg_out [7:0];
  assign _107_ = \aes_reg_key0_i.en ? aes_key0_dataout : 8'b00000000;
  assign _108_ = \aes_reg_ctr_i.en ? aes_ctr_dataout : _107_;
  assign _109_ = \aes_reg_oplen_i.en ? aes_len_dataout : _108_;
  assign _110_ = \aes_reg_opaddr_i.en ? aes_addr_dataout : _109_;
  logic [7:0] fangyuan0;
  assign fangyuan0 = { 6'b000000, aes_reg_state };
  assign data_out = sel_reg_state ? fangyuan0 : _110_;
  assign _014_[15:0] = _033_ ? _008_ : operated_bytes_count;
  assign operated_bytes_count_next = reset_byte_counter ? 16'b0000000000000000 : _014_[15:0];
  assign _111_[15:0] = more_blocks ? _009_ : block_counter;
  assign block_counter_next = reset_byte_counter ? 16'b0000000000000000 : _111_[15:0];
  assign _112_[3:0] = xram_ack ? _010_ : byte_counter;
  assign byte_counter_next = reset_byte_counter ? 4'b0000 : _112_[3:0];
  assign aes_reg_state_next_read_data = last_byte_acked ? 2'b10 : 2'b01;
  assign _113_ = last_byte_acked ? 2'b00 : 2'b11;
  assign aes_reg_state_next_write_data = _034_ ? 2'b01 : _113_;
  assign _114_ = aes_state_write_data ? aes_reg_state_next_write_data : 2'b00;
  logic [1:0] fangyuan1;
  assign fangyuan1 = { 1'b1, aes_time_enough };
  assign _115_ = aes_state_operate ? fangyuan1 : _114_;
  assign _116_ = aes_state_read_data ? aes_reg_state_next_read_data : _115_;
  logic [1:0] fangyuan2;
  assign fangyuan2 = { 1'b0, reset_byte_counter };
  assign aes_reg_state_next = aes_state_idle ? fangyuan2 : _116_;
  assign mem_data_buf_next[7:0] = _035_ ? xram_data_in : mem_data_buf[7:0];
  assign mem_data_buf_next[15:8] = _036_ ? xram_data_in : mem_data_buf[15:8];
  assign mem_data_buf_next[23:16] = _037_ ? xram_data_in : mem_data_buf[23:16];
  assign mem_data_buf_next[31:24] = _038_ ? xram_data_in : mem_data_buf[31:24];
  assign mem_data_buf_next[39:32] = _039_ ? xram_data_in : mem_data_buf[39:32];
  assign mem_data_buf_next[47:40] = _040_ ? xram_data_in : mem_data_buf[47:40];
  assign mem_data_buf_next[55:48] = _041_ ? xram_data_in : mem_data_buf[55:48];
  assign mem_data_buf_next[63:56] = _042_ ? xram_data_in : mem_data_buf[63:56];
  assign mem_data_buf_next[71:64] = _043_ ? xram_data_in : mem_data_buf[71:64];
  assign mem_data_buf_next[79:72] = _044_ ? xram_data_in : mem_data_buf[79:72];
  assign mem_data_buf_next[87:80] = _045_ ? xram_data_in : mem_data_buf[87:80];
  assign mem_data_buf_next[95:88] = _046_ ? xram_data_in : mem_data_buf[95:88];
  assign mem_data_buf_next[103:96] = _047_ ? xram_data_in : mem_data_buf[103:96];
  assign mem_data_buf_next[111:104] = _048_ ? xram_data_in : mem_data_buf[111:104];
  assign mem_data_buf_next[119:112] = _049_ ? xram_data_in : mem_data_buf[119:112];
  assign mem_data_buf_next[127:120] = last_byte_acked ? xram_data_in : mem_data_buf[127:120];
  assign _117_ = more_blocks ? _012_ : uaes_ctr;
  assign uaes_ctr_nxt = reset_byte_counter ? \aes_reg_ctr_i.reg_out : _117_;
  assign _118_ = _053_ ? _013_ : aes_time_counter;
  assign aes_time_counter_next = _050_ ? 5'b00000 : _118_;
  assign encrypted_data_buf_next = aes_state_operate ? encrypted_data : encrypted_data_buf;
  assign _119_ = _030_ ? encrypted_data_buf[119:112] : encrypted_data_buf[127:120];
  assign _120_ = _029_ ? encrypted_data_buf[111:104] : _119_;
  assign _121_ = _028_ ? encrypted_data_buf[103:96] : _120_;
  assign _122_ = _027_ ? encrypted_data_buf[95:88] : _121_;
  assign _123_ = _026_ ? encrypted_data_buf[87:80] : _122_;
  assign _124_ = _025_ ? encrypted_data_buf[79:72] : _123_;
  assign _125_ = _024_ ? encrypted_data_buf[71:64] : _124_;
  assign _126_ = _023_ ? encrypted_data_buf[63:56] : _125_;
  assign _127_ = _022_ ? encrypted_data_buf[55:48] : _126_;
  assign _128_ = _021_ ? encrypted_data_buf[47:40] : _127_;
  assign _129_ = _020_ ? encrypted_data_buf[39:32] : _128_;
  assign _130_ = _019_ ? encrypted_data_buf[31:24] : _129_;
  assign _131_ = _018_ ? encrypted_data_buf[23:16] : _130_;
  assign _132_ = _017_ ? encrypted_data_buf[15:8] : _131_;
  assign xram_data_out = _016_ ? encrypted_data_buf[7:0] : _132_;
  assign encrypted_data = aes_out ^ mem_data_buf;
  aes_128 aes_128_i (
    .clk(clk),
    .key(\aes_reg_key0_i.reg_out ),
    .out(aes_out),
    .state(uaes_ctr)
  );
  assign aes_addr = \aes_reg_opaddr_i.reg_out ;
  assign aes_ctr = \aes_reg_ctr_i.reg_out ;
  assign aes_curr_key = \aes_reg_key0_i.reg_out ;
  assign aes_key0 = \aes_reg_key0_i.reg_out ;
  assign aes_len = \aes_reg_oplen_i.reg_out ;
  assign aes_reg_ctr = \aes_reg_ctr_i.reg_out ;
  assign \aes_reg_ctr_i.addr = addr[3:0];
  assign \aes_reg_ctr_i.clk = clk;
  assign \aes_reg_ctr_i.data_in = data_in;
  assign \aes_reg_ctr_i.data_out = aes_ctr_dataout;
  assign \aes_reg_ctr_i.data_out_mux = aes_ctr_dataout;
  assign \aes_reg_ctr_i.rst = rst;
  assign aes_reg_key0 = \aes_reg_key0_i.reg_out ;
  assign \aes_reg_key0_i.addr = addr[3:0];
  assign \aes_reg_key0_i.clk = clk;
  assign \aes_reg_key0_i.data_in = data_in;
  assign \aes_reg_key0_i.data_out = aes_key0_dataout;
  assign \aes_reg_key0_i.data_out_mux = aes_key0_dataout;
  assign \aes_reg_key0_i.rst = rst;
  assign aes_reg_opaddr = \aes_reg_opaddr_i.reg_out ;
  assign \aes_reg_opaddr_i.addr = addr[0];
  assign \aes_reg_opaddr_i.clk = clk;
  assign \aes_reg_opaddr_i.data_in = data_in;
  assign \aes_reg_opaddr_i.data_out = aes_addr_dataout;
  assign \aes_reg_opaddr_i.data_out_mux = aes_addr_dataout;
  assign \aes_reg_opaddr_i.rst = rst;
  assign aes_reg_oplen = \aes_reg_oplen_i.reg_out ;
  assign \aes_reg_oplen_i.addr = addr[0];
  assign \aes_reg_oplen_i.clk = clk;
  assign \aes_reg_oplen_i.data_in = data_in;
  assign \aes_reg_oplen_i.data_out = aes_len_dataout;
  assign \aes_reg_oplen_i.data_out_mux = aes_len_dataout;
  assign \aes_reg_oplen_i.rst = rst;
  assign aes_reg_state_next_idle = reset_byte_counter;
  assign aes_reg_state_next_operate = aes_time_enough;
  assign aes_state = aes_reg_state;
  assign incr_byte_counter = xram_ack;
  assign sel_reg_addr = \aes_reg_opaddr_i.en ;
  assign sel_reg_ctr = \aes_reg_ctr_i.en ;
  assign sel_reg_key0 = \aes_reg_key0_i.en ;
  assign sel_reg_len = \aes_reg_oplen_i.en ;
  assign start_op = reset_byte_counter;
  assign xram_wr = aes_state_write_data;
endmodule
