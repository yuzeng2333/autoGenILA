module SDP_X_chn_trt_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:2129" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:2130" *)
  output outsig;
  assign outsig = in_0;
endmodule
