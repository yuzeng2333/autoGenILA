module NV_BLKBOX_SRC0(Y);
  (* src = "/u/yuzeng/nvdla1/hw/outdir/nv_full/vmod/vlibs/NV_BLKBOX_SRC0.v:12" *)
  output Y;
  assign Y = 1'b0;
  assign Y = Y ~^ Y;
endmodule
