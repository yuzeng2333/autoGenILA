module FP17_TO_FP32_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_to_fp32.v:85" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp32.v:86" *)
  output outsig;
  assign outsig = in_0;
endmodule
