module NV_NVDLA_CMAC_CORE_rt_in(nvdla_core_clk, nvdla_core_rstn, sc2mac_dat_data0, sc2mac_dat_data1, sc2mac_dat_data10, sc2mac_dat_data100, sc2mac_dat_data101, sc2mac_dat_data102, sc2mac_dat_data103, sc2mac_dat_data104, sc2mac_dat_data105, sc2mac_dat_data106, sc2mac_dat_data107, sc2mac_dat_data108, sc2mac_dat_data109, sc2mac_dat_data11, sc2mac_dat_data110, sc2mac_dat_data111, sc2mac_dat_data112, sc2mac_dat_data113, sc2mac_dat_data114, sc2mac_dat_data115, sc2mac_dat_data116, sc2mac_dat_data117, sc2mac_dat_data118, sc2mac_dat_data119, sc2mac_dat_data12, sc2mac_dat_data120, sc2mac_dat_data121, sc2mac_dat_data122, sc2mac_dat_data123, sc2mac_dat_data124, sc2mac_dat_data125, sc2mac_dat_data126, sc2mac_dat_data127, sc2mac_dat_data13, sc2mac_dat_data14, sc2mac_dat_data15, sc2mac_dat_data16, sc2mac_dat_data17, sc2mac_dat_data18, sc2mac_dat_data19, sc2mac_dat_data2, sc2mac_dat_data20, sc2mac_dat_data21, sc2mac_dat_data22, sc2mac_dat_data23, sc2mac_dat_data24, sc2mac_dat_data25, sc2mac_dat_data26, sc2mac_dat_data27, sc2mac_dat_data28, sc2mac_dat_data29, sc2mac_dat_data3, sc2mac_dat_data30, sc2mac_dat_data31, sc2mac_dat_data32, sc2mac_dat_data33, sc2mac_dat_data34, sc2mac_dat_data35, sc2mac_dat_data36, sc2mac_dat_data37, sc2mac_dat_data38, sc2mac_dat_data39, sc2mac_dat_data4, sc2mac_dat_data40, sc2mac_dat_data41, sc2mac_dat_data42, sc2mac_dat_data43, sc2mac_dat_data44, sc2mac_dat_data45, sc2mac_dat_data46, sc2mac_dat_data47, sc2mac_dat_data48, sc2mac_dat_data49, sc2mac_dat_data5, sc2mac_dat_data50, sc2mac_dat_data51, sc2mac_dat_data52, sc2mac_dat_data53, sc2mac_dat_data54, sc2mac_dat_data55, sc2mac_dat_data56, sc2mac_dat_data57, sc2mac_dat_data58, sc2mac_dat_data59, sc2mac_dat_data6, sc2mac_dat_data60, sc2mac_dat_data61, sc2mac_dat_data62, sc2mac_dat_data63, sc2mac_dat_data64, sc2mac_dat_data65, sc2mac_dat_data66, sc2mac_dat_data67, sc2mac_dat_data68, sc2mac_dat_data69, sc2mac_dat_data7, sc2mac_dat_data70, sc2mac_dat_data71, sc2mac_dat_data72, sc2mac_dat_data73, sc2mac_dat_data74, sc2mac_dat_data75, sc2mac_dat_data76, sc2mac_dat_data77, sc2mac_dat_data78, sc2mac_dat_data79, sc2mac_dat_data8, sc2mac_dat_data80, sc2mac_dat_data81, sc2mac_dat_data82, sc2mac_dat_data83, sc2mac_dat_data84, sc2mac_dat_data85, sc2mac_dat_data86, sc2mac_dat_data87, sc2mac_dat_data88, sc2mac_dat_data89, sc2mac_dat_data9, sc2mac_dat_data90, sc2mac_dat_data91, sc2mac_dat_data92, sc2mac_dat_data93, sc2mac_dat_data94, sc2mac_dat_data95, sc2mac_dat_data96, sc2mac_dat_data97, sc2mac_dat_data98, sc2mac_dat_data99, sc2mac_dat_mask, sc2mac_dat_pd, sc2mac_dat_pvld, sc2mac_wt_data0, sc2mac_wt_data1, sc2mac_wt_data10, sc2mac_wt_data100, sc2mac_wt_data101, sc2mac_wt_data102, sc2mac_wt_data103, sc2mac_wt_data104, sc2mac_wt_data105, sc2mac_wt_data106, sc2mac_wt_data107, sc2mac_wt_data108, sc2mac_wt_data109, sc2mac_wt_data11, sc2mac_wt_data110, sc2mac_wt_data111, sc2mac_wt_data112, sc2mac_wt_data113, sc2mac_wt_data114, sc2mac_wt_data115, sc2mac_wt_data116, sc2mac_wt_data117, sc2mac_wt_data118, sc2mac_wt_data119, sc2mac_wt_data12, sc2mac_wt_data120, sc2mac_wt_data121, sc2mac_wt_data122, sc2mac_wt_data123, sc2mac_wt_data124, sc2mac_wt_data125, sc2mac_wt_data126, sc2mac_wt_data127, sc2mac_wt_data13, sc2mac_wt_data14, sc2mac_wt_data15, sc2mac_wt_data16, sc2mac_wt_data17, sc2mac_wt_data18, sc2mac_wt_data19, sc2mac_wt_data2, sc2mac_wt_data20, sc2mac_wt_data21, sc2mac_wt_data22, sc2mac_wt_data23, sc2mac_wt_data24, sc2mac_wt_data25, sc2mac_wt_data26, sc2mac_wt_data27, sc2mac_wt_data28, sc2mac_wt_data29, sc2mac_wt_data3, sc2mac_wt_data30, sc2mac_wt_data31, sc2mac_wt_data32, sc2mac_wt_data33, sc2mac_wt_data34, sc2mac_wt_data35, sc2mac_wt_data36, sc2mac_wt_data37, sc2mac_wt_data38, sc2mac_wt_data39, sc2mac_wt_data4, sc2mac_wt_data40, sc2mac_wt_data41, sc2mac_wt_data42, sc2mac_wt_data43, sc2mac_wt_data44, sc2mac_wt_data45, sc2mac_wt_data46, sc2mac_wt_data47, sc2mac_wt_data48, sc2mac_wt_data49, sc2mac_wt_data5, sc2mac_wt_data50, sc2mac_wt_data51, sc2mac_wt_data52, sc2mac_wt_data53, sc2mac_wt_data54, sc2mac_wt_data55, sc2mac_wt_data56, sc2mac_wt_data57, sc2mac_wt_data58, sc2mac_wt_data59, sc2mac_wt_data6, sc2mac_wt_data60, sc2mac_wt_data61, sc2mac_wt_data62, sc2mac_wt_data63, sc2mac_wt_data64, sc2mac_wt_data65, sc2mac_wt_data66, sc2mac_wt_data67, sc2mac_wt_data68, sc2mac_wt_data69, sc2mac_wt_data7, sc2mac_wt_data70, sc2mac_wt_data71, sc2mac_wt_data72, sc2mac_wt_data73, sc2mac_wt_data74, sc2mac_wt_data75, sc2mac_wt_data76, sc2mac_wt_data77, sc2mac_wt_data78, sc2mac_wt_data79, sc2mac_wt_data8, sc2mac_wt_data80, sc2mac_wt_data81, sc2mac_wt_data82, sc2mac_wt_data83, sc2mac_wt_data84, sc2mac_wt_data85, sc2mac_wt_data86, sc2mac_wt_data87, sc2mac_wt_data88, sc2mac_wt_data89, sc2mac_wt_data9, sc2mac_wt_data90, sc2mac_wt_data91, sc2mac_wt_data92, sc2mac_wt_data93, sc2mac_wt_data94, sc2mac_wt_data95, sc2mac_wt_data96, sc2mac_wt_data97, sc2mac_wt_data98, sc2mac_wt_data99, sc2mac_wt_mask, sc2mac_wt_pvld, sc2mac_wt_sel, in_dat_data0, in_dat_data1, in_dat_data10, in_dat_data100, in_dat_data101, in_dat_data102, in_dat_data103, in_dat_data104, in_dat_data105, in_dat_data106, in_dat_data107, in_dat_data108, in_dat_data109, in_dat_data11, in_dat_data110, in_dat_data111, in_dat_data112, in_dat_data113, in_dat_data114, in_dat_data115, in_dat_data116, in_dat_data117, in_dat_data118, in_dat_data119, in_dat_data12, in_dat_data120, in_dat_data121, in_dat_data122, in_dat_data123, in_dat_data124, in_dat_data125, in_dat_data126, in_dat_data127, in_dat_data13, in_dat_data14, in_dat_data15, in_dat_data16, in_dat_data17, in_dat_data18, in_dat_data19, in_dat_data2, in_dat_data20, in_dat_data21, in_dat_data22, in_dat_data23, in_dat_data24, in_dat_data25, in_dat_data26, in_dat_data27, in_dat_data28, in_dat_data29, in_dat_data3, in_dat_data30, in_dat_data31, in_dat_data32, in_dat_data33, in_dat_data34, in_dat_data35, in_dat_data36, in_dat_data37, in_dat_data38, in_dat_data39, in_dat_data4, in_dat_data40, in_dat_data41, in_dat_data42, in_dat_data43, in_dat_data44, in_dat_data45, in_dat_data46, in_dat_data47, in_dat_data48, in_dat_data49, in_dat_data5, in_dat_data50, in_dat_data51, in_dat_data52, in_dat_data53, in_dat_data54, in_dat_data55, in_dat_data56, in_dat_data57, in_dat_data58, in_dat_data59, in_dat_data6, in_dat_data60, in_dat_data61, in_dat_data62, in_dat_data63, in_dat_data64, in_dat_data65, in_dat_data66, in_dat_data67, in_dat_data68, in_dat_data69, in_dat_data7, in_dat_data70, in_dat_data71, in_dat_data72, in_dat_data73, in_dat_data74, in_dat_data75, in_dat_data76, in_dat_data77, in_dat_data78, in_dat_data79, in_dat_data8, in_dat_data80, in_dat_data81, in_dat_data82, in_dat_data83, in_dat_data84, in_dat_data85, in_dat_data86, in_dat_data87, in_dat_data88, in_dat_data89, in_dat_data9, in_dat_data90, in_dat_data91, in_dat_data92, in_dat_data93, in_dat_data94, in_dat_data95, in_dat_data96, in_dat_data97, in_dat_data98, in_dat_data99, in_dat_mask, in_dat_pd, in_dat_pvld, in_dat_stripe_end, in_dat_stripe_st, in_wt_data0, in_wt_data1, in_wt_data10, in_wt_data100, in_wt_data101, in_wt_data102, in_wt_data103, in_wt_data104, in_wt_data105, in_wt_data106, in_wt_data107, in_wt_data108, in_wt_data109, in_wt_data11, in_wt_data110, in_wt_data111, in_wt_data112, in_wt_data113, in_wt_data114, in_wt_data115, in_wt_data116, in_wt_data117, in_wt_data118, in_wt_data119, in_wt_data12, in_wt_data120, in_wt_data121, in_wt_data122, in_wt_data123, in_wt_data124, in_wt_data125, in_wt_data126, in_wt_data127, in_wt_data13, in_wt_data14, in_wt_data15, in_wt_data16, in_wt_data17, in_wt_data18, in_wt_data19, in_wt_data2, in_wt_data20, in_wt_data21, in_wt_data22, in_wt_data23, in_wt_data24, in_wt_data25, in_wt_data26, in_wt_data27, in_wt_data28, in_wt_data29, in_wt_data3, in_wt_data30, in_wt_data31, in_wt_data32, in_wt_data33, in_wt_data34, in_wt_data35, in_wt_data36, in_wt_data37, in_wt_data38, in_wt_data39, in_wt_data4, in_wt_data40, in_wt_data41, in_wt_data42, in_wt_data43, in_wt_data44, in_wt_data45, in_wt_data46, in_wt_data47, in_wt_data48, in_wt_data49, in_wt_data5, in_wt_data50, in_wt_data51, in_wt_data52, in_wt_data53, in_wt_data54, in_wt_data55, in_wt_data56, in_wt_data57, in_wt_data58, in_wt_data59, in_wt_data6, in_wt_data60, in_wt_data61, in_wt_data62, in_wt_data63, in_wt_data64, in_wt_data65, in_wt_data66, in_wt_data67, in_wt_data68, in_wt_data69, in_wt_data7, in_wt_data70, in_wt_data71, in_wt_data72, in_wt_data73, in_wt_data74, in_wt_data75, in_wt_data76, in_wt_data77, in_wt_data78, in_wt_data79, in_wt_data8, in_wt_data80, in_wt_data81, in_wt_data82, in_wt_data83, in_wt_data84, in_wt_data85, in_wt_data86, in_wt_data87, in_wt_data88, in_wt_data89, in_wt_data9, in_wt_data90, in_wt_data91, in_wt_data92, in_wt_data93, in_wt_data94, in_wt_data95, in_wt_data96, in_wt_data97, in_wt_data98, in_wt_data99, in_wt_mask, in_wt_pvld, in_wt_sel);
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3018" *)
  wire [7:0] _000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3028" *)
  wire [7:0] _001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3038" *)
  wire [7:0] _002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1888" *)
  wire [7:0] _003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1898" *)
  wire [7:0] _004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1908" *)
  wire [7:0] _005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1918" *)
  wire [7:0] _006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1928" *)
  wire [7:0] _007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1938" *)
  wire [7:0] _008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1948" *)
  wire [7:0] _009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1958" *)
  wire [7:0] _010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1778" *)
  wire [7:0] _011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1968" *)
  wire [7:0] _012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1978" *)
  wire [7:0] _013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1988" *)
  wire [7:0] _014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1998" *)
  wire [7:0] _015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2008" *)
  wire [7:0] _016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2018" *)
  wire [7:0] _017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2028" *)
  wire [7:0] _018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2038" *)
  wire [7:0] _019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2048" *)
  wire [7:0] _020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2058" *)
  wire [7:0] _021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1788" *)
  wire [7:0] _022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2068" *)
  wire [7:0] _023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2078" *)
  wire [7:0] _024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2088" *)
  wire [7:0] _025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2098" *)
  wire [7:0] _026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2108" *)
  wire [7:0] _027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2118" *)
  wire [7:0] _028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2128" *)
  wire [7:0] _029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2138" *)
  wire [7:0] _030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2148" *)
  wire [7:0] _031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2158" *)
  wire [7:0] _032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1798" *)
  wire [7:0] _033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2168" *)
  wire [7:0] _034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2178" *)
  wire [7:0] _035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2188" *)
  wire [7:0] _036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2198" *)
  wire [7:0] _037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2208" *)
  wire [7:0] _038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2218" *)
  wire [7:0] _039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2228" *)
  wire [7:0] _040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2238" *)
  wire [7:0] _041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2248" *)
  wire [7:0] _042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2258" *)
  wire [7:0] _043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1808" *)
  wire [7:0] _044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2268" *)
  wire [7:0] _045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2278" *)
  wire [7:0] _046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2288" *)
  wire [7:0] _047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2298" *)
  wire [7:0] _048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2308" *)
  wire [7:0] _049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2318" *)
  wire [7:0] _050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2328" *)
  wire [7:0] _051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2338" *)
  wire [7:0] _052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2348" *)
  wire [7:0] _053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2358" *)
  wire [7:0] _054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1818" *)
  wire [7:0] _055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2368" *)
  wire [7:0] _056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2378" *)
  wire [7:0] _057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2388" *)
  wire [7:0] _058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2398" *)
  wire [7:0] _059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2408" *)
  wire [7:0] _060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2418" *)
  wire [7:0] _061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2428" *)
  wire [7:0] _062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2438" *)
  wire [7:0] _063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2448" *)
  wire [7:0] _064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2458" *)
  wire [7:0] _065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1828" *)
  wire [7:0] _066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2468" *)
  wire [7:0] _067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2478" *)
  wire [7:0] _068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2488" *)
  wire [7:0] _069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2498" *)
  wire [7:0] _070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2508" *)
  wire [7:0] _071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2518" *)
  wire [7:0] _072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2528" *)
  wire [7:0] _073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2538" *)
  wire [7:0] _074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2548" *)
  wire [7:0] _075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2558" *)
  wire [7:0] _076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1838" *)
  wire [7:0] _077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2568" *)
  wire [7:0] _078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2578" *)
  wire [7:0] _079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2588" *)
  wire [7:0] _080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2598" *)
  wire [7:0] _081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2608" *)
  wire [7:0] _082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2618" *)
  wire [7:0] _083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2628" *)
  wire [7:0] _084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2638" *)
  wire [7:0] _085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2648" *)
  wire [7:0] _086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2658" *)
  wire [7:0] _087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1848" *)
  wire [7:0] _088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2668" *)
  wire [7:0] _089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2678" *)
  wire [7:0] _090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2688" *)
  wire [7:0] _091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2698" *)
  wire [7:0] _092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2708" *)
  wire [7:0] _093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2718" *)
  wire [7:0] _094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2728" *)
  wire [7:0] _095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2738" *)
  wire [7:0] _096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2748" *)
  wire [7:0] _097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2758" *)
  wire [7:0] _098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1858" *)
  wire [7:0] _099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1768" *)
  wire [7:0] _100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2768" *)
  wire [7:0] _101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2778" *)
  wire [7:0] _102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2788" *)
  wire [7:0] _103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2798" *)
  wire [7:0] _104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2808" *)
  wire [7:0] _105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2818" *)
  wire [7:0] _106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2828" *)
  wire [7:0] _107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2838" *)
  wire [7:0] _108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2848" *)
  wire [7:0] _109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2858" *)
  wire [7:0] _110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1868" *)
  wire [7:0] _111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2868" *)
  wire [7:0] _112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2878" *)
  wire [7:0] _113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2888" *)
  wire [7:0] _114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2898" *)
  wire [7:0] _115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2908" *)
  wire [7:0] _116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2918" *)
  wire [7:0] _117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2928" *)
  wire [7:0] _118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2938" *)
  wire [7:0] _119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2948" *)
  wire [7:0] _120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2958" *)
  wire [7:0] _121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1878" *)
  wire [7:0] _122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2968" *)
  wire [7:0] _123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2978" *)
  wire [7:0] _124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2988" *)
  wire [7:0] _125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2998" *)
  wire [7:0] _126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3008" *)
  wire [7:0] _127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1646" *)
  wire [127:0] _128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1707" *)
  wire [8:0] _129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4427" *)
  wire [7:0] _130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4437" *)
  wire [7:0] _131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4447" *)
  wire [7:0] _132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3297" *)
  wire [7:0] _133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3307" *)
  wire [7:0] _134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3317" *)
  wire [7:0] _135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3327" *)
  wire [7:0] _136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3337" *)
  wire [7:0] _137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3347" *)
  wire [7:0] _138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3357" *)
  wire [7:0] _139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3367" *)
  wire [7:0] _140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3187" *)
  wire [7:0] _141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3377" *)
  wire [7:0] _142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3387" *)
  wire [7:0] _143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3397" *)
  wire [7:0] _144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3407" *)
  wire [7:0] _145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3417" *)
  wire [7:0] _146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3427" *)
  wire [7:0] _147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3437" *)
  wire [7:0] _148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3447" *)
  wire [7:0] _149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3457" *)
  wire [7:0] _150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3467" *)
  wire [7:0] _151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3197" *)
  wire [7:0] _152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3477" *)
  wire [7:0] _153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3487" *)
  wire [7:0] _154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3497" *)
  wire [7:0] _155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3507" *)
  wire [7:0] _156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3517" *)
  wire [7:0] _157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3527" *)
  wire [7:0] _158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3537" *)
  wire [7:0] _159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3547" *)
  wire [7:0] _160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3557" *)
  wire [7:0] _161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3567" *)
  wire [7:0] _162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3207" *)
  wire [7:0] _163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3577" *)
  wire [7:0] _164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3587" *)
  wire [7:0] _165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3597" *)
  wire [7:0] _166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3607" *)
  wire [7:0] _167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3617" *)
  wire [7:0] _168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3627" *)
  wire [7:0] _169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3637" *)
  wire [7:0] _170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3647" *)
  wire [7:0] _171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3657" *)
  wire [7:0] _172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3667" *)
  wire [7:0] _173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3217" *)
  wire [7:0] _174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3677" *)
  wire [7:0] _175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3687" *)
  wire [7:0] _176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3697" *)
  wire [7:0] _177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3707" *)
  wire [7:0] _178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3717" *)
  wire [7:0] _179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3727" *)
  wire [7:0] _180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3737" *)
  wire [7:0] _181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3747" *)
  wire [7:0] _182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3757" *)
  wire [7:0] _183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3767" *)
  wire [7:0] _184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3227" *)
  wire [7:0] _185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3777" *)
  wire [7:0] _186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3787" *)
  wire [7:0] _187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3797" *)
  wire [7:0] _188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3807" *)
  wire [7:0] _189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3817" *)
  wire [7:0] _190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3827" *)
  wire [7:0] _191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3837" *)
  wire [7:0] _192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3847" *)
  wire [7:0] _193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3857" *)
  wire [7:0] _194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3867" *)
  wire [7:0] _195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3237" *)
  wire [7:0] _196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3877" *)
  wire [7:0] _197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3887" *)
  wire [7:0] _198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3897" *)
  wire [7:0] _199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3907" *)
  wire [7:0] _200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3917" *)
  wire [7:0] _201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3927" *)
  wire [7:0] _202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3937" *)
  wire [7:0] _203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3947" *)
  wire [7:0] _204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3957" *)
  wire [7:0] _205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3967" *)
  wire [7:0] _206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3247" *)
  wire [7:0] _207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3977" *)
  wire [7:0] _208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3987" *)
  wire [7:0] _209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3997" *)
  wire [7:0] _210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4007" *)
  wire [7:0] _211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4017" *)
  wire [7:0] _212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4027" *)
  wire [7:0] _213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4037" *)
  wire [7:0] _214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4047" *)
  wire [7:0] _215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4057" *)
  wire [7:0] _216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4067" *)
  wire [7:0] _217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3257" *)
  wire [7:0] _218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4077" *)
  wire [7:0] _219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4087" *)
  wire [7:0] _220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4097" *)
  wire [7:0] _221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4107" *)
  wire [7:0] _222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4117" *)
  wire [7:0] _223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4127" *)
  wire [7:0] _224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4137" *)
  wire [7:0] _225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4147" *)
  wire [7:0] _226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4157" *)
  wire [7:0] _227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4167" *)
  wire [7:0] _228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3267" *)
  wire [7:0] _229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3177" *)
  wire [7:0] _230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4177" *)
  wire [7:0] _231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4187" *)
  wire [7:0] _232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4197" *)
  wire [7:0] _233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4207" *)
  wire [7:0] _234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4217" *)
  wire [7:0] _235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4227" *)
  wire [7:0] _236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4237" *)
  wire [7:0] _237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4247" *)
  wire [7:0] _238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4257" *)
  wire [7:0] _239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4267" *)
  wire [7:0] _240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3277" *)
  wire [7:0] _241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4277" *)
  wire [7:0] _242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4287" *)
  wire [7:0] _243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4297" *)
  wire [7:0] _244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4307" *)
  wire [7:0] _245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4317" *)
  wire [7:0] _246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4327" *)
  wire [7:0] _247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4337" *)
  wire [7:0] _248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4347" *)
  wire [7:0] _249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4357" *)
  wire [7:0] _250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4367" *)
  wire [7:0] _251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3287" *)
  wire [7:0] _252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4377" *)
  wire [7:0] _253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4387" *)
  wire [7:0] _254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4397" *)
  wire [7:0] _255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4407" *)
  wire [7:0] _256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4417" *)
  wire [7:0] _257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3116" *)
  wire [127:0] _258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3055" *)
  wire [7:0] _259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1650" *)
  wire _260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3059" *)
  wire _261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1067" *)
  wire [1023:0] in_dat_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:803" *)
  output [7:0] in_dat_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:804" *)
  output [7:0] in_dat_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:805" *)
  output [7:0] in_dat_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:806" *)
  output [7:0] in_dat_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:807" *)
  output [7:0] in_dat_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:808" *)
  output [7:0] in_dat_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:809" *)
  output [7:0] in_dat_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:810" *)
  output [7:0] in_dat_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:811" *)
  output [7:0] in_dat_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:812" *)
  output [7:0] in_dat_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:813" *)
  output [7:0] in_dat_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:814" *)
  output [7:0] in_dat_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:815" *)
  output [7:0] in_dat_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:816" *)
  output [7:0] in_dat_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:817" *)
  output [7:0] in_dat_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:818" *)
  output [7:0] in_dat_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:819" *)
  output [7:0] in_dat_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:820" *)
  output [7:0] in_dat_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:821" *)
  output [7:0] in_dat_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:822" *)
  output [7:0] in_dat_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:823" *)
  output [7:0] in_dat_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:824" *)
  output [7:0] in_dat_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:825" *)
  output [7:0] in_dat_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:826" *)
  output [7:0] in_dat_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:827" *)
  output [7:0] in_dat_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:828" *)
  output [7:0] in_dat_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:829" *)
  output [7:0] in_dat_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:830" *)
  output [7:0] in_dat_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:831" *)
  output [7:0] in_dat_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:832" *)
  output [7:0] in_dat_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:833" *)
  output [7:0] in_dat_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:834" *)
  output [7:0] in_dat_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:835" *)
  output [7:0] in_dat_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:836" *)
  output [7:0] in_dat_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:837" *)
  output [7:0] in_dat_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:838" *)
  output [7:0] in_dat_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:839" *)
  output [7:0] in_dat_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:840" *)
  output [7:0] in_dat_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:841" *)
  output [7:0] in_dat_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:842" *)
  output [7:0] in_dat_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:843" *)
  output [7:0] in_dat_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:844" *)
  output [7:0] in_dat_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:845" *)
  output [7:0] in_dat_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:846" *)
  output [7:0] in_dat_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:847" *)
  output [7:0] in_dat_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:848" *)
  output [7:0] in_dat_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:849" *)
  output [7:0] in_dat_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:850" *)
  output [7:0] in_dat_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:851" *)
  output [7:0] in_dat_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:852" *)
  output [7:0] in_dat_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:853" *)
  output [7:0] in_dat_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:854" *)
  output [7:0] in_dat_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:855" *)
  output [7:0] in_dat_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:856" *)
  output [7:0] in_dat_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:857" *)
  output [7:0] in_dat_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:858" *)
  output [7:0] in_dat_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:859" *)
  output [7:0] in_dat_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:860" *)
  output [7:0] in_dat_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:861" *)
  output [7:0] in_dat_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:862" *)
  output [7:0] in_dat_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:863" *)
  output [7:0] in_dat_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:864" *)
  output [7:0] in_dat_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:865" *)
  output [7:0] in_dat_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:866" *)
  output [7:0] in_dat_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:867" *)
  output [7:0] in_dat_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:868" *)
  output [7:0] in_dat_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:869" *)
  output [7:0] in_dat_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:870" *)
  output [7:0] in_dat_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:871" *)
  output [7:0] in_dat_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:872" *)
  output [7:0] in_dat_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:873" *)
  output [7:0] in_dat_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:874" *)
  output [7:0] in_dat_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:875" *)
  output [7:0] in_dat_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:876" *)
  output [7:0] in_dat_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:877" *)
  output [7:0] in_dat_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:878" *)
  output [7:0] in_dat_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:879" *)
  output [7:0] in_dat_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:880" *)
  output [7:0] in_dat_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:881" *)
  output [7:0] in_dat_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:882" *)
  output [7:0] in_dat_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:883" *)
  output [7:0] in_dat_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:884" *)
  output [7:0] in_dat_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:885" *)
  output [7:0] in_dat_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:886" *)
  output [7:0] in_dat_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:887" *)
  output [7:0] in_dat_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:888" *)
  output [7:0] in_dat_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:889" *)
  output [7:0] in_dat_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:890" *)
  output [7:0] in_dat_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:891" *)
  output [7:0] in_dat_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:892" *)
  output [7:0] in_dat_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:893" *)
  output [7:0] in_dat_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:894" *)
  output [7:0] in_dat_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:895" *)
  output [7:0] in_dat_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:896" *)
  output [7:0] in_dat_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:897" *)
  output [7:0] in_dat_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:898" *)
  output [7:0] in_dat_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:899" *)
  output [7:0] in_dat_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:900" *)
  output [7:0] in_dat_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:901" *)
  output [7:0] in_dat_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:902" *)
  output [7:0] in_dat_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:903" *)
  output [7:0] in_dat_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:904" *)
  output [7:0] in_dat_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:905" *)
  output [7:0] in_dat_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:906" *)
  output [7:0] in_dat_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:907" *)
  output [7:0] in_dat_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:908" *)
  output [7:0] in_dat_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:909" *)
  output [7:0] in_dat_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:910" *)
  output [7:0] in_dat_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:911" *)
  output [7:0] in_dat_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:912" *)
  output [7:0] in_dat_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:913" *)
  output [7:0] in_dat_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:914" *)
  output [7:0] in_dat_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:915" *)
  output [7:0] in_dat_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:916" *)
  output [7:0] in_dat_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:917" *)
  output [7:0] in_dat_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:918" *)
  output [7:0] in_dat_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:919" *)
  output [7:0] in_dat_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:920" *)
  output [7:0] in_dat_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:921" *)
  output [7:0] in_dat_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:922" *)
  output [7:0] in_dat_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:923" *)
  output [7:0] in_dat_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:924" *)
  output [7:0] in_dat_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:925" *)
  output [7:0] in_dat_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:926" *)
  output [7:0] in_dat_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:927" *)
  output [7:0] in_dat_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:928" *)
  output [7:0] in_dat_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:929" *)
  output [7:0] in_dat_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:930" *)
  output [7:0] in_dat_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:931" *)
  output [127:0] in_dat_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:932" *)
  output [8:0] in_dat_pd;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:933" *)
  output in_dat_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:934" *)
  output in_dat_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:935" *)
  output in_dat_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1201" *)
  wire [1023:0] in_rt_dat_data_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1202" *)
  reg [1023:0] in_rt_dat_data_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1203" *)
  wire [127:0] in_rt_dat_mask_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1204" *)
  reg [127:0] in_rt_dat_mask_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1205" *)
  wire [8:0] in_rt_dat_pd_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1206" *)
  reg [8:0] in_rt_dat_pd_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1207" *)
  wire in_rt_dat_pvld_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1208" *)
  reg in_rt_dat_pvld_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1209" *)
  wire [1023:0] in_rt_wt_data_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1210" *)
  reg [1023:0] in_rt_wt_data_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1211" *)
  wire [127:0] in_rt_wt_mask_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1212" *)
  reg [127:0] in_rt_wt_mask_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1213" *)
  wire in_rt_wt_pvld_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1214" *)
  reg in_rt_wt_pvld_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1215" *)
  wire [7:0] in_rt_wt_sel_d0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1216" *)
  reg [7:0] in_rt_wt_sel_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1217" *)
  wire [1023:0] in_wt_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:936" *)
  output [7:0] in_wt_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:937" *)
  output [7:0] in_wt_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:938" *)
  output [7:0] in_wt_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:939" *)
  output [7:0] in_wt_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:940" *)
  output [7:0] in_wt_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:941" *)
  output [7:0] in_wt_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:942" *)
  output [7:0] in_wt_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:943" *)
  output [7:0] in_wt_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:944" *)
  output [7:0] in_wt_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:945" *)
  output [7:0] in_wt_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:946" *)
  output [7:0] in_wt_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:947" *)
  output [7:0] in_wt_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:948" *)
  output [7:0] in_wt_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:949" *)
  output [7:0] in_wt_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:950" *)
  output [7:0] in_wt_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:951" *)
  output [7:0] in_wt_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:952" *)
  output [7:0] in_wt_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:953" *)
  output [7:0] in_wt_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:954" *)
  output [7:0] in_wt_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:955" *)
  output [7:0] in_wt_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:956" *)
  output [7:0] in_wt_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:957" *)
  output [7:0] in_wt_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:958" *)
  output [7:0] in_wt_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:959" *)
  output [7:0] in_wt_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:960" *)
  output [7:0] in_wt_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:961" *)
  output [7:0] in_wt_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:962" *)
  output [7:0] in_wt_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:963" *)
  output [7:0] in_wt_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:964" *)
  output [7:0] in_wt_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:965" *)
  output [7:0] in_wt_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:966" *)
  output [7:0] in_wt_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:967" *)
  output [7:0] in_wt_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:968" *)
  output [7:0] in_wt_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:969" *)
  output [7:0] in_wt_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:970" *)
  output [7:0] in_wt_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:971" *)
  output [7:0] in_wt_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:972" *)
  output [7:0] in_wt_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:973" *)
  output [7:0] in_wt_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:974" *)
  output [7:0] in_wt_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:975" *)
  output [7:0] in_wt_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:976" *)
  output [7:0] in_wt_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:977" *)
  output [7:0] in_wt_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:978" *)
  output [7:0] in_wt_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:979" *)
  output [7:0] in_wt_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:980" *)
  output [7:0] in_wt_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:981" *)
  output [7:0] in_wt_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:982" *)
  output [7:0] in_wt_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:983" *)
  output [7:0] in_wt_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:984" *)
  output [7:0] in_wt_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:985" *)
  output [7:0] in_wt_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:986" *)
  output [7:0] in_wt_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:987" *)
  output [7:0] in_wt_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:988" *)
  output [7:0] in_wt_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:989" *)
  output [7:0] in_wt_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:990" *)
  output [7:0] in_wt_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:991" *)
  output [7:0] in_wt_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:992" *)
  output [7:0] in_wt_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:993" *)
  output [7:0] in_wt_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:994" *)
  output [7:0] in_wt_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:995" *)
  output [7:0] in_wt_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:996" *)
  output [7:0] in_wt_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:997" *)
  output [7:0] in_wt_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:998" *)
  output [7:0] in_wt_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:999" *)
  output [7:0] in_wt_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1000" *)
  output [7:0] in_wt_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1001" *)
  output [7:0] in_wt_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1002" *)
  output [7:0] in_wt_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1003" *)
  output [7:0] in_wt_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1004" *)
  output [7:0] in_wt_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1005" *)
  output [7:0] in_wt_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1006" *)
  output [7:0] in_wt_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1007" *)
  output [7:0] in_wt_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1008" *)
  output [7:0] in_wt_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1009" *)
  output [7:0] in_wt_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1010" *)
  output [7:0] in_wt_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1011" *)
  output [7:0] in_wt_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1012" *)
  output [7:0] in_wt_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1013" *)
  output [7:0] in_wt_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1014" *)
  output [7:0] in_wt_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1015" *)
  output [7:0] in_wt_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1016" *)
  output [7:0] in_wt_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1017" *)
  output [7:0] in_wt_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1018" *)
  output [7:0] in_wt_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1019" *)
  output [7:0] in_wt_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1020" *)
  output [7:0] in_wt_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1021" *)
  output [7:0] in_wt_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1022" *)
  output [7:0] in_wt_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1023" *)
  output [7:0] in_wt_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1024" *)
  output [7:0] in_wt_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1025" *)
  output [7:0] in_wt_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1026" *)
  output [7:0] in_wt_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1027" *)
  output [7:0] in_wt_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1028" *)
  output [7:0] in_wt_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1029" *)
  output [7:0] in_wt_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1030" *)
  output [7:0] in_wt_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1031" *)
  output [7:0] in_wt_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1032" *)
  output [7:0] in_wt_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1033" *)
  output [7:0] in_wt_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1034" *)
  output [7:0] in_wt_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1035" *)
  output [7:0] in_wt_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1036" *)
  output [7:0] in_wt_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1037" *)
  output [7:0] in_wt_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1038" *)
  output [7:0] in_wt_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1039" *)
  output [7:0] in_wt_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1040" *)
  output [7:0] in_wt_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1041" *)
  output [7:0] in_wt_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1042" *)
  output [7:0] in_wt_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1043" *)
  output [7:0] in_wt_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1044" *)
  output [7:0] in_wt_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1045" *)
  output [7:0] in_wt_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1046" *)
  output [7:0] in_wt_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1047" *)
  output [7:0] in_wt_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1048" *)
  output [7:0] in_wt_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1049" *)
  output [7:0] in_wt_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1050" *)
  output [7:0] in_wt_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1051" *)
  output [7:0] in_wt_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1052" *)
  output [7:0] in_wt_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1053" *)
  output [7:0] in_wt_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1054" *)
  output [7:0] in_wt_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1055" *)
  output [7:0] in_wt_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1056" *)
  output [7:0] in_wt_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1057" *)
  output [7:0] in_wt_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1058" *)
  output [7:0] in_wt_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1059" *)
  output [7:0] in_wt_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1060" *)
  output [7:0] in_wt_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1061" *)
  output [7:0] in_wt_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1062" *)
  output [7:0] in_wt_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1063" *)
  output [7:0] in_wt_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1064" *)
  output [127:0] in_wt_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1065" *)
  output in_wt_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1066" *)
  output [7:0] in_wt_sel;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:539" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:540" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:541" *)
  input [7:0] sc2mac_dat_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:542" *)
  input [7:0] sc2mac_dat_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:543" *)
  input [7:0] sc2mac_dat_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:544" *)
  input [7:0] sc2mac_dat_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:545" *)
  input [7:0] sc2mac_dat_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:546" *)
  input [7:0] sc2mac_dat_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:547" *)
  input [7:0] sc2mac_dat_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:548" *)
  input [7:0] sc2mac_dat_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:549" *)
  input [7:0] sc2mac_dat_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:550" *)
  input [7:0] sc2mac_dat_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:551" *)
  input [7:0] sc2mac_dat_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:552" *)
  input [7:0] sc2mac_dat_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:553" *)
  input [7:0] sc2mac_dat_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:554" *)
  input [7:0] sc2mac_dat_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:555" *)
  input [7:0] sc2mac_dat_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:556" *)
  input [7:0] sc2mac_dat_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:557" *)
  input [7:0] sc2mac_dat_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:558" *)
  input [7:0] sc2mac_dat_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:559" *)
  input [7:0] sc2mac_dat_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:560" *)
  input [7:0] sc2mac_dat_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:561" *)
  input [7:0] sc2mac_dat_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:562" *)
  input [7:0] sc2mac_dat_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:563" *)
  input [7:0] sc2mac_dat_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:564" *)
  input [7:0] sc2mac_dat_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:565" *)
  input [7:0] sc2mac_dat_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:566" *)
  input [7:0] sc2mac_dat_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:567" *)
  input [7:0] sc2mac_dat_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:568" *)
  input [7:0] sc2mac_dat_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:569" *)
  input [7:0] sc2mac_dat_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:570" *)
  input [7:0] sc2mac_dat_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:571" *)
  input [7:0] sc2mac_dat_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:572" *)
  input [7:0] sc2mac_dat_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:573" *)
  input [7:0] sc2mac_dat_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:574" *)
  input [7:0] sc2mac_dat_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:575" *)
  input [7:0] sc2mac_dat_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:576" *)
  input [7:0] sc2mac_dat_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:577" *)
  input [7:0] sc2mac_dat_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:578" *)
  input [7:0] sc2mac_dat_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:579" *)
  input [7:0] sc2mac_dat_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:580" *)
  input [7:0] sc2mac_dat_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:581" *)
  input [7:0] sc2mac_dat_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:582" *)
  input [7:0] sc2mac_dat_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:583" *)
  input [7:0] sc2mac_dat_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:584" *)
  input [7:0] sc2mac_dat_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:585" *)
  input [7:0] sc2mac_dat_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:586" *)
  input [7:0] sc2mac_dat_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:587" *)
  input [7:0] sc2mac_dat_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:588" *)
  input [7:0] sc2mac_dat_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:589" *)
  input [7:0] sc2mac_dat_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:590" *)
  input [7:0] sc2mac_dat_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:591" *)
  input [7:0] sc2mac_dat_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:592" *)
  input [7:0] sc2mac_dat_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:593" *)
  input [7:0] sc2mac_dat_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:594" *)
  input [7:0] sc2mac_dat_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:595" *)
  input [7:0] sc2mac_dat_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:596" *)
  input [7:0] sc2mac_dat_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:597" *)
  input [7:0] sc2mac_dat_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:598" *)
  input [7:0] sc2mac_dat_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:599" *)
  input [7:0] sc2mac_dat_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:600" *)
  input [7:0] sc2mac_dat_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:601" *)
  input [7:0] sc2mac_dat_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:602" *)
  input [7:0] sc2mac_dat_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:603" *)
  input [7:0] sc2mac_dat_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:604" *)
  input [7:0] sc2mac_dat_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:605" *)
  input [7:0] sc2mac_dat_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:606" *)
  input [7:0] sc2mac_dat_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:607" *)
  input [7:0] sc2mac_dat_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:608" *)
  input [7:0] sc2mac_dat_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:609" *)
  input [7:0] sc2mac_dat_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:610" *)
  input [7:0] sc2mac_dat_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:611" *)
  input [7:0] sc2mac_dat_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:612" *)
  input [7:0] sc2mac_dat_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:613" *)
  input [7:0] sc2mac_dat_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:614" *)
  input [7:0] sc2mac_dat_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:615" *)
  input [7:0] sc2mac_dat_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:616" *)
  input [7:0] sc2mac_dat_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:617" *)
  input [7:0] sc2mac_dat_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:618" *)
  input [7:0] sc2mac_dat_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:619" *)
  input [7:0] sc2mac_dat_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:620" *)
  input [7:0] sc2mac_dat_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:621" *)
  input [7:0] sc2mac_dat_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:622" *)
  input [7:0] sc2mac_dat_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:623" *)
  input [7:0] sc2mac_dat_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:624" *)
  input [7:0] sc2mac_dat_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:625" *)
  input [7:0] sc2mac_dat_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:626" *)
  input [7:0] sc2mac_dat_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:627" *)
  input [7:0] sc2mac_dat_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:628" *)
  input [7:0] sc2mac_dat_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:629" *)
  input [7:0] sc2mac_dat_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:630" *)
  input [7:0] sc2mac_dat_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:631" *)
  input [7:0] sc2mac_dat_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:632" *)
  input [7:0] sc2mac_dat_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:633" *)
  input [7:0] sc2mac_dat_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:634" *)
  input [7:0] sc2mac_dat_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:635" *)
  input [7:0] sc2mac_dat_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:636" *)
  input [7:0] sc2mac_dat_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:637" *)
  input [7:0] sc2mac_dat_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:638" *)
  input [7:0] sc2mac_dat_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:639" *)
  input [7:0] sc2mac_dat_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:640" *)
  input [7:0] sc2mac_dat_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:641" *)
  input [7:0] sc2mac_dat_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:642" *)
  input [7:0] sc2mac_dat_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:643" *)
  input [7:0] sc2mac_dat_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:644" *)
  input [7:0] sc2mac_dat_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:645" *)
  input [7:0] sc2mac_dat_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:646" *)
  input [7:0] sc2mac_dat_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:647" *)
  input [7:0] sc2mac_dat_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:648" *)
  input [7:0] sc2mac_dat_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:649" *)
  input [7:0] sc2mac_dat_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:650" *)
  input [7:0] sc2mac_dat_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:651" *)
  input [7:0] sc2mac_dat_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:652" *)
  input [7:0] sc2mac_dat_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:653" *)
  input [7:0] sc2mac_dat_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:654" *)
  input [7:0] sc2mac_dat_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:655" *)
  input [7:0] sc2mac_dat_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:656" *)
  input [7:0] sc2mac_dat_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:657" *)
  input [7:0] sc2mac_dat_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:658" *)
  input [7:0] sc2mac_dat_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:659" *)
  input [7:0] sc2mac_dat_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:660" *)
  input [7:0] sc2mac_dat_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:661" *)
  input [7:0] sc2mac_dat_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:662" *)
  input [7:0] sc2mac_dat_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:663" *)
  input [7:0] sc2mac_dat_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:664" *)
  input [7:0] sc2mac_dat_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:665" *)
  input [7:0] sc2mac_dat_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:666" *)
  input [7:0] sc2mac_dat_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:667" *)
  input [7:0] sc2mac_dat_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:668" *)
  input [7:0] sc2mac_dat_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:669" *)
  input [127:0] sc2mac_dat_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:670" *)
  input [8:0] sc2mac_dat_pd;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:671" *)
  input sc2mac_dat_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:672" *)
  input [7:0] sc2mac_wt_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:673" *)
  input [7:0] sc2mac_wt_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:674" *)
  input [7:0] sc2mac_wt_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:675" *)
  input [7:0] sc2mac_wt_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:676" *)
  input [7:0] sc2mac_wt_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:677" *)
  input [7:0] sc2mac_wt_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:678" *)
  input [7:0] sc2mac_wt_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:679" *)
  input [7:0] sc2mac_wt_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:680" *)
  input [7:0] sc2mac_wt_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:681" *)
  input [7:0] sc2mac_wt_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:682" *)
  input [7:0] sc2mac_wt_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:683" *)
  input [7:0] sc2mac_wt_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:684" *)
  input [7:0] sc2mac_wt_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:685" *)
  input [7:0] sc2mac_wt_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:686" *)
  input [7:0] sc2mac_wt_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:687" *)
  input [7:0] sc2mac_wt_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:688" *)
  input [7:0] sc2mac_wt_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:689" *)
  input [7:0] sc2mac_wt_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:690" *)
  input [7:0] sc2mac_wt_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:691" *)
  input [7:0] sc2mac_wt_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:692" *)
  input [7:0] sc2mac_wt_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:693" *)
  input [7:0] sc2mac_wt_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:694" *)
  input [7:0] sc2mac_wt_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:695" *)
  input [7:0] sc2mac_wt_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:696" *)
  input [7:0] sc2mac_wt_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:697" *)
  input [7:0] sc2mac_wt_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:698" *)
  input [7:0] sc2mac_wt_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:699" *)
  input [7:0] sc2mac_wt_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:700" *)
  input [7:0] sc2mac_wt_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:701" *)
  input [7:0] sc2mac_wt_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:702" *)
  input [7:0] sc2mac_wt_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:703" *)
  input [7:0] sc2mac_wt_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:704" *)
  input [7:0] sc2mac_wt_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:705" *)
  input [7:0] sc2mac_wt_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:706" *)
  input [7:0] sc2mac_wt_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:707" *)
  input [7:0] sc2mac_wt_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:708" *)
  input [7:0] sc2mac_wt_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:709" *)
  input [7:0] sc2mac_wt_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:710" *)
  input [7:0] sc2mac_wt_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:711" *)
  input [7:0] sc2mac_wt_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:712" *)
  input [7:0] sc2mac_wt_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:713" *)
  input [7:0] sc2mac_wt_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:714" *)
  input [7:0] sc2mac_wt_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:715" *)
  input [7:0] sc2mac_wt_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:716" *)
  input [7:0] sc2mac_wt_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:717" *)
  input [7:0] sc2mac_wt_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:718" *)
  input [7:0] sc2mac_wt_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:719" *)
  input [7:0] sc2mac_wt_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:720" *)
  input [7:0] sc2mac_wt_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:721" *)
  input [7:0] sc2mac_wt_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:722" *)
  input [7:0] sc2mac_wt_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:723" *)
  input [7:0] sc2mac_wt_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:724" *)
  input [7:0] sc2mac_wt_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:725" *)
  input [7:0] sc2mac_wt_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:726" *)
  input [7:0] sc2mac_wt_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:727" *)
  input [7:0] sc2mac_wt_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:728" *)
  input [7:0] sc2mac_wt_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:729" *)
  input [7:0] sc2mac_wt_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:730" *)
  input [7:0] sc2mac_wt_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:731" *)
  input [7:0] sc2mac_wt_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:732" *)
  input [7:0] sc2mac_wt_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:733" *)
  input [7:0] sc2mac_wt_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:734" *)
  input [7:0] sc2mac_wt_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:735" *)
  input [7:0] sc2mac_wt_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:736" *)
  input [7:0] sc2mac_wt_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:737" *)
  input [7:0] sc2mac_wt_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:738" *)
  input [7:0] sc2mac_wt_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:739" *)
  input [7:0] sc2mac_wt_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:740" *)
  input [7:0] sc2mac_wt_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:741" *)
  input [7:0] sc2mac_wt_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:742" *)
  input [7:0] sc2mac_wt_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:743" *)
  input [7:0] sc2mac_wt_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:744" *)
  input [7:0] sc2mac_wt_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:745" *)
  input [7:0] sc2mac_wt_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:746" *)
  input [7:0] sc2mac_wt_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:747" *)
  input [7:0] sc2mac_wt_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:748" *)
  input [7:0] sc2mac_wt_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:749" *)
  input [7:0] sc2mac_wt_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:750" *)
  input [7:0] sc2mac_wt_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:751" *)
  input [7:0] sc2mac_wt_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:752" *)
  input [7:0] sc2mac_wt_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:753" *)
  input [7:0] sc2mac_wt_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:754" *)
  input [7:0] sc2mac_wt_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:755" *)
  input [7:0] sc2mac_wt_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:756" *)
  input [7:0] sc2mac_wt_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:757" *)
  input [7:0] sc2mac_wt_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:758" *)
  input [7:0] sc2mac_wt_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:759" *)
  input [7:0] sc2mac_wt_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:760" *)
  input [7:0] sc2mac_wt_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:761" *)
  input [7:0] sc2mac_wt_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:762" *)
  input [7:0] sc2mac_wt_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:763" *)
  input [7:0] sc2mac_wt_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:764" *)
  input [7:0] sc2mac_wt_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:765" *)
  input [7:0] sc2mac_wt_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:766" *)
  input [7:0] sc2mac_wt_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:767" *)
  input [7:0] sc2mac_wt_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:768" *)
  input [7:0] sc2mac_wt_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:769" *)
  input [7:0] sc2mac_wt_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:770" *)
  input [7:0] sc2mac_wt_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:771" *)
  input [7:0] sc2mac_wt_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:772" *)
  input [7:0] sc2mac_wt_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:773" *)
  input [7:0] sc2mac_wt_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:774" *)
  input [7:0] sc2mac_wt_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:775" *)
  input [7:0] sc2mac_wt_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:776" *)
  input [7:0] sc2mac_wt_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:777" *)
  input [7:0] sc2mac_wt_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:778" *)
  input [7:0] sc2mac_wt_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:779" *)
  input [7:0] sc2mac_wt_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:780" *)
  input [7:0] sc2mac_wt_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:781" *)
  input [7:0] sc2mac_wt_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:782" *)
  input [7:0] sc2mac_wt_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:783" *)
  input [7:0] sc2mac_wt_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:784" *)
  input [7:0] sc2mac_wt_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:785" *)
  input [7:0] sc2mac_wt_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:786" *)
  input [7:0] sc2mac_wt_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:787" *)
  input [7:0] sc2mac_wt_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:788" *)
  input [7:0] sc2mac_wt_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:789" *)
  input [7:0] sc2mac_wt_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:790" *)
  input [7:0] sc2mac_wt_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:791" *)
  input [7:0] sc2mac_wt_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:792" *)
  input [7:0] sc2mac_wt_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:793" *)
  input [7:0] sc2mac_wt_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:794" *)
  input [7:0] sc2mac_wt_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:795" *)
  input [7:0] sc2mac_wt_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:796" *)
  input [7:0] sc2mac_wt_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:797" *)
  input [7:0] sc2mac_wt_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:798" *)
  input [7:0] sc2mac_wt_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:799" *)
  input [7:0] sc2mac_wt_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:800" *)
  input [127:0] sc2mac_wt_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:801" *)
  input sc2mac_wt_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:802" *)
  input [7:0] sc2mac_wt_sel;
  assign _260_ = sc2mac_dat_pvld | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1650" *) in_rt_dat_pvld_d1;
  assign _261_ = sc2mac_wt_pvld | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3059" *) in_rt_wt_pvld_d1;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[1023:1016] <= _132_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[1015:1008] <= _131_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[1007:1000] <= _130_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[999:992] <= _257_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[991:984] <= _256_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[983:976] <= _255_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[975:968] <= _254_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[967:960] <= _253_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[959:952] <= _251_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[951:944] <= _250_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[943:936] <= _249_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[935:928] <= _248_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[927:920] <= _247_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[919:912] <= _246_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[911:904] <= _245_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[903:896] <= _244_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[895:888] <= _243_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[887:880] <= _242_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[879:872] <= _240_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[871:864] <= _239_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[863:856] <= _238_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[855:848] <= _237_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[847:840] <= _236_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[839:832] <= _235_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[831:824] <= _234_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[823:816] <= _233_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[815:808] <= _232_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[807:800] <= _231_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[799:792] <= _228_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[791:784] <= _227_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[783:776] <= _226_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[775:768] <= _225_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[767:760] <= _224_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[759:752] <= _223_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[751:744] <= _222_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[743:736] <= _221_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[735:728] <= _220_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[727:720] <= _219_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[719:712] <= _217_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[711:704] <= _216_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[703:696] <= _215_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[695:688] <= _214_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[687:680] <= _213_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[679:672] <= _212_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[671:664] <= _211_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[663:656] <= _210_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[655:648] <= _209_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[647:640] <= _208_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[639:632] <= _206_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[631:624] <= _205_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[623:616] <= _204_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[615:608] <= _203_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[607:600] <= _202_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[599:592] <= _201_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[591:584] <= _200_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[583:576] <= _199_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[575:568] <= _198_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[567:560] <= _197_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[559:552] <= _195_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[551:544] <= _194_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[543:536] <= _193_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[535:528] <= _192_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[527:520] <= _191_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[519:512] <= _190_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[511:504] <= _189_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[503:496] <= _188_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[495:488] <= _187_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[487:480] <= _186_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[479:472] <= _184_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[471:464] <= _183_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[463:456] <= _182_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[455:448] <= _181_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[447:440] <= _180_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[439:432] <= _179_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[431:424] <= _178_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[423:416] <= _177_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[415:408] <= _176_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[407:400] <= _175_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[399:392] <= _173_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[391:384] <= _172_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[383:376] <= _171_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[375:368] <= _170_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[367:360] <= _169_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[359:352] <= _168_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[351:344] <= _167_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[343:336] <= _166_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[335:328] <= _165_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[327:320] <= _164_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[319:312] <= _162_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[311:304] <= _161_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[303:296] <= _160_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[295:288] <= _159_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[287:280] <= _158_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[279:272] <= _157_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[271:264] <= _156_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[263:256] <= _155_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[255:248] <= _154_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[247:240] <= _153_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[239:232] <= _151_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[231:224] <= _150_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[223:216] <= _149_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[215:208] <= _148_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[207:200] <= _147_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[199:192] <= _146_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[191:184] <= _145_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[183:176] <= _144_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[175:168] <= _143_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[167:160] <= _142_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[159:152] <= _140_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[151:144] <= _139_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[143:136] <= _138_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[135:128] <= _137_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[127:120] <= _136_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[119:112] <= _135_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[111:104] <= _134_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[103:96] <= _133_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[95:88] <= _252_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[87:80] <= _241_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[79:72] <= _229_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[71:64] <= _218_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[63:56] <= _207_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[55:48] <= _196_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[47:40] <= _185_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[39:32] <= _174_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[31:24] <= _163_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[23:16] <= _152_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[15:8] <= _141_;
  always @(posedge nvdla_core_clk)
      in_rt_wt_data_d1[7:0] <= _230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_wt_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      in_rt_wt_mask_d1 <= _258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_wt_sel_d1 <= 8'b00000000;
    else
      in_rt_wt_sel_d1 <= _259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_wt_pvld_d1 <= 1'b0;
    else
      in_rt_wt_pvld_d1 <= sc2mac_wt_pvld;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[1023:1016] <= _002_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[1015:1008] <= _001_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[1007:1000] <= _000_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[999:992] <= _127_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[991:984] <= _126_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[983:976] <= _125_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[975:968] <= _124_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[967:960] <= _123_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[959:952] <= _121_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[951:944] <= _120_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[943:936] <= _119_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[935:928] <= _118_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[927:920] <= _117_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[919:912] <= _116_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[911:904] <= _115_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[903:896] <= _114_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[895:888] <= _113_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[887:880] <= _112_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[879:872] <= _110_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[871:864] <= _109_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[863:856] <= _108_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[855:848] <= _107_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[847:840] <= _106_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[839:832] <= _105_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[831:824] <= _104_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[823:816] <= _103_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[815:808] <= _102_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[807:800] <= _101_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[799:792] <= _098_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[791:784] <= _097_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[783:776] <= _096_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[775:768] <= _095_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[767:760] <= _094_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[759:752] <= _093_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[751:744] <= _092_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[743:736] <= _091_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[735:728] <= _090_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[727:720] <= _089_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[719:712] <= _087_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[711:704] <= _086_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[703:696] <= _085_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[695:688] <= _084_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[687:680] <= _083_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[679:672] <= _082_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[671:664] <= _081_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[663:656] <= _080_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[655:648] <= _079_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[647:640] <= _078_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[639:632] <= _076_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[631:624] <= _075_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[623:616] <= _074_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[615:608] <= _073_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[607:600] <= _072_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[599:592] <= _071_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[591:584] <= _070_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[583:576] <= _069_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[575:568] <= _068_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[567:560] <= _067_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[559:552] <= _065_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[551:544] <= _064_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[543:536] <= _063_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[535:528] <= _062_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[527:520] <= _061_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[519:512] <= _060_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[511:504] <= _059_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[503:496] <= _058_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[495:488] <= _057_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[487:480] <= _056_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[479:472] <= _054_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[471:464] <= _053_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[463:456] <= _052_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[455:448] <= _051_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[447:440] <= _050_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[439:432] <= _049_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[431:424] <= _048_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[423:416] <= _047_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[415:408] <= _046_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[407:400] <= _045_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[399:392] <= _043_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[391:384] <= _042_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[383:376] <= _041_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[375:368] <= _040_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[367:360] <= _039_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[359:352] <= _038_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[351:344] <= _037_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[343:336] <= _036_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[335:328] <= _035_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[327:320] <= _034_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[319:312] <= _032_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[311:304] <= _031_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[303:296] <= _030_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[295:288] <= _029_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[287:280] <= _028_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[279:272] <= _027_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[271:264] <= _026_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[263:256] <= _025_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[255:248] <= _024_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[247:240] <= _023_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[239:232] <= _021_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[231:224] <= _020_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[223:216] <= _019_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[215:208] <= _018_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[207:200] <= _017_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[199:192] <= _016_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[191:184] <= _015_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[183:176] <= _014_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[175:168] <= _013_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[167:160] <= _012_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[159:152] <= _010_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[151:144] <= _009_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[143:136] <= _008_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[135:128] <= _007_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[127:120] <= _006_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[119:112] <= _005_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[111:104] <= _004_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[103:96] <= _003_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[95:88] <= _122_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[87:80] <= _111_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[79:72] <= _099_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[71:64] <= _088_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[63:56] <= _077_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[55:48] <= _066_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[47:40] <= _055_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[39:32] <= _044_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[31:24] <= _033_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[23:16] <= _022_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[15:8] <= _011_;
  always @(posedge nvdla_core_clk)
      in_rt_dat_data_d1[7:0] <= _100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_dat_pd_d1 <= 9'b000000000;
    else
      in_rt_dat_pd_d1 <= _129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_dat_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      in_rt_dat_mask_d1 <= _128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      in_rt_dat_pvld_d1 <= 1'b0;
    else
      in_rt_dat_pvld_d1 <= sc2mac_dat_pvld;
  assign _132_ = sc2mac_wt_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4448" *) sc2mac_wt_data127 : in_rt_wt_data_d1[1023:1016];
  assign _131_ = sc2mac_wt_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4438" *) sc2mac_wt_data126 : in_rt_wt_data_d1[1015:1008];
  assign _130_ = sc2mac_wt_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4428" *) sc2mac_wt_data125 : in_rt_wt_data_d1[1007:1000];
  assign _257_ = sc2mac_wt_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4418" *) sc2mac_wt_data124 : in_rt_wt_data_d1[999:992];
  assign _256_ = sc2mac_wt_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4408" *) sc2mac_wt_data123 : in_rt_wt_data_d1[991:984];
  assign _255_ = sc2mac_wt_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4398" *) sc2mac_wt_data122 : in_rt_wt_data_d1[983:976];
  assign _254_ = sc2mac_wt_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4388" *) sc2mac_wt_data121 : in_rt_wt_data_d1[975:968];
  assign _253_ = sc2mac_wt_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4378" *) sc2mac_wt_data120 : in_rt_wt_data_d1[967:960];
  assign _251_ = sc2mac_wt_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4368" *) sc2mac_wt_data119 : in_rt_wt_data_d1[959:952];
  assign _250_ = sc2mac_wt_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4358" *) sc2mac_wt_data118 : in_rt_wt_data_d1[951:944];
  assign _249_ = sc2mac_wt_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4348" *) sc2mac_wt_data117 : in_rt_wt_data_d1[943:936];
  assign _248_ = sc2mac_wt_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4338" *) sc2mac_wt_data116 : in_rt_wt_data_d1[935:928];
  assign _247_ = sc2mac_wt_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4328" *) sc2mac_wt_data115 : in_rt_wt_data_d1[927:920];
  assign _246_ = sc2mac_wt_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4318" *) sc2mac_wt_data114 : in_rt_wt_data_d1[919:912];
  assign _245_ = sc2mac_wt_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4308" *) sc2mac_wt_data113 : in_rt_wt_data_d1[911:904];
  assign _244_ = sc2mac_wt_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4298" *) sc2mac_wt_data112 : in_rt_wt_data_d1[903:896];
  assign _243_ = sc2mac_wt_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4288" *) sc2mac_wt_data111 : in_rt_wt_data_d1[895:888];
  assign _242_ = sc2mac_wt_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4278" *) sc2mac_wt_data110 : in_rt_wt_data_d1[887:880];
  assign _240_ = sc2mac_wt_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4268" *) sc2mac_wt_data109 : in_rt_wt_data_d1[879:872];
  assign _239_ = sc2mac_wt_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4258" *) sc2mac_wt_data108 : in_rt_wt_data_d1[871:864];
  assign _238_ = sc2mac_wt_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4248" *) sc2mac_wt_data107 : in_rt_wt_data_d1[863:856];
  assign _237_ = sc2mac_wt_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4238" *) sc2mac_wt_data106 : in_rt_wt_data_d1[855:848];
  assign _236_ = sc2mac_wt_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4228" *) sc2mac_wt_data105 : in_rt_wt_data_d1[847:840];
  assign _235_ = sc2mac_wt_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4218" *) sc2mac_wt_data104 : in_rt_wt_data_d1[839:832];
  assign _234_ = sc2mac_wt_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4208" *) sc2mac_wt_data103 : in_rt_wt_data_d1[831:824];
  assign _233_ = sc2mac_wt_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4198" *) sc2mac_wt_data102 : in_rt_wt_data_d1[823:816];
  assign _232_ = sc2mac_wt_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4188" *) sc2mac_wt_data101 : in_rt_wt_data_d1[815:808];
  assign _231_ = sc2mac_wt_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4178" *) sc2mac_wt_data100 : in_rt_wt_data_d1[807:800];
  assign _228_ = sc2mac_wt_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4168" *) sc2mac_wt_data99 : in_rt_wt_data_d1[799:792];
  assign _227_ = sc2mac_wt_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4158" *) sc2mac_wt_data98 : in_rt_wt_data_d1[791:784];
  assign _226_ = sc2mac_wt_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4148" *) sc2mac_wt_data97 : in_rt_wt_data_d1[783:776];
  assign _225_ = sc2mac_wt_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4138" *) sc2mac_wt_data96 : in_rt_wt_data_d1[775:768];
  assign _224_ = sc2mac_wt_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4128" *) sc2mac_wt_data95 : in_rt_wt_data_d1[767:760];
  assign _223_ = sc2mac_wt_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4118" *) sc2mac_wt_data94 : in_rt_wt_data_d1[759:752];
  assign _222_ = sc2mac_wt_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4108" *) sc2mac_wt_data93 : in_rt_wt_data_d1[751:744];
  assign _221_ = sc2mac_wt_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4098" *) sc2mac_wt_data92 : in_rt_wt_data_d1[743:736];
  assign _220_ = sc2mac_wt_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4088" *) sc2mac_wt_data91 : in_rt_wt_data_d1[735:728];
  assign _219_ = sc2mac_wt_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4078" *) sc2mac_wt_data90 : in_rt_wt_data_d1[727:720];
  assign _217_ = sc2mac_wt_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4068" *) sc2mac_wt_data89 : in_rt_wt_data_d1[719:712];
  assign _216_ = sc2mac_wt_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4058" *) sc2mac_wt_data88 : in_rt_wt_data_d1[711:704];
  assign _215_ = sc2mac_wt_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4048" *) sc2mac_wt_data87 : in_rt_wt_data_d1[703:696];
  assign _214_ = sc2mac_wt_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4038" *) sc2mac_wt_data86 : in_rt_wt_data_d1[695:688];
  assign _213_ = sc2mac_wt_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4028" *) sc2mac_wt_data85 : in_rt_wt_data_d1[687:680];
  assign _212_ = sc2mac_wt_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4018" *) sc2mac_wt_data84 : in_rt_wt_data_d1[679:672];
  assign _211_ = sc2mac_wt_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:4008" *) sc2mac_wt_data83 : in_rt_wt_data_d1[671:664];
  assign _210_ = sc2mac_wt_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3998" *) sc2mac_wt_data82 : in_rt_wt_data_d1[663:656];
  assign _209_ = sc2mac_wt_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3988" *) sc2mac_wt_data81 : in_rt_wt_data_d1[655:648];
  assign _208_ = sc2mac_wt_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3978" *) sc2mac_wt_data80 : in_rt_wt_data_d1[647:640];
  assign _206_ = sc2mac_wt_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3968" *) sc2mac_wt_data79 : in_rt_wt_data_d1[639:632];
  assign _205_ = sc2mac_wt_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3958" *) sc2mac_wt_data78 : in_rt_wt_data_d1[631:624];
  assign _204_ = sc2mac_wt_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3948" *) sc2mac_wt_data77 : in_rt_wt_data_d1[623:616];
  assign _203_ = sc2mac_wt_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3938" *) sc2mac_wt_data76 : in_rt_wt_data_d1[615:608];
  assign _202_ = sc2mac_wt_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3928" *) sc2mac_wt_data75 : in_rt_wt_data_d1[607:600];
  assign _201_ = sc2mac_wt_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3918" *) sc2mac_wt_data74 : in_rt_wt_data_d1[599:592];
  assign _200_ = sc2mac_wt_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3908" *) sc2mac_wt_data73 : in_rt_wt_data_d1[591:584];
  assign _199_ = sc2mac_wt_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3898" *) sc2mac_wt_data72 : in_rt_wt_data_d1[583:576];
  assign _198_ = sc2mac_wt_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3888" *) sc2mac_wt_data71 : in_rt_wt_data_d1[575:568];
  assign _197_ = sc2mac_wt_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3878" *) sc2mac_wt_data70 : in_rt_wt_data_d1[567:560];
  assign _195_ = sc2mac_wt_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3868" *) sc2mac_wt_data69 : in_rt_wt_data_d1[559:552];
  assign _194_ = sc2mac_wt_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3858" *) sc2mac_wt_data68 : in_rt_wt_data_d1[551:544];
  assign _193_ = sc2mac_wt_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3848" *) sc2mac_wt_data67 : in_rt_wt_data_d1[543:536];
  assign _192_ = sc2mac_wt_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3838" *) sc2mac_wt_data66 : in_rt_wt_data_d1[535:528];
  assign _191_ = sc2mac_wt_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3828" *) sc2mac_wt_data65 : in_rt_wt_data_d1[527:520];
  assign _190_ = sc2mac_wt_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3818" *) sc2mac_wt_data64 : in_rt_wt_data_d1[519:512];
  assign _189_ = sc2mac_wt_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3808" *) sc2mac_wt_data63 : in_rt_wt_data_d1[511:504];
  assign _188_ = sc2mac_wt_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3798" *) sc2mac_wt_data62 : in_rt_wt_data_d1[503:496];
  assign _187_ = sc2mac_wt_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3788" *) sc2mac_wt_data61 : in_rt_wt_data_d1[495:488];
  assign _186_ = sc2mac_wt_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3778" *) sc2mac_wt_data60 : in_rt_wt_data_d1[487:480];
  assign _184_ = sc2mac_wt_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3768" *) sc2mac_wt_data59 : in_rt_wt_data_d1[479:472];
  assign _183_ = sc2mac_wt_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3758" *) sc2mac_wt_data58 : in_rt_wt_data_d1[471:464];
  assign _182_ = sc2mac_wt_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3748" *) sc2mac_wt_data57 : in_rt_wt_data_d1[463:456];
  assign _181_ = sc2mac_wt_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3738" *) sc2mac_wt_data56 : in_rt_wt_data_d1[455:448];
  assign _180_ = sc2mac_wt_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3728" *) sc2mac_wt_data55 : in_rt_wt_data_d1[447:440];
  assign _179_ = sc2mac_wt_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3718" *) sc2mac_wt_data54 : in_rt_wt_data_d1[439:432];
  assign _178_ = sc2mac_wt_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3708" *) sc2mac_wt_data53 : in_rt_wt_data_d1[431:424];
  assign _177_ = sc2mac_wt_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3698" *) sc2mac_wt_data52 : in_rt_wt_data_d1[423:416];
  assign _176_ = sc2mac_wt_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3688" *) sc2mac_wt_data51 : in_rt_wt_data_d1[415:408];
  assign _175_ = sc2mac_wt_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3678" *) sc2mac_wt_data50 : in_rt_wt_data_d1[407:400];
  assign _173_ = sc2mac_wt_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3668" *) sc2mac_wt_data49 : in_rt_wt_data_d1[399:392];
  assign _172_ = sc2mac_wt_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3658" *) sc2mac_wt_data48 : in_rt_wt_data_d1[391:384];
  assign _171_ = sc2mac_wt_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3648" *) sc2mac_wt_data47 : in_rt_wt_data_d1[383:376];
  assign _170_ = sc2mac_wt_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3638" *) sc2mac_wt_data46 : in_rt_wt_data_d1[375:368];
  assign _169_ = sc2mac_wt_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3628" *) sc2mac_wt_data45 : in_rt_wt_data_d1[367:360];
  assign _168_ = sc2mac_wt_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3618" *) sc2mac_wt_data44 : in_rt_wt_data_d1[359:352];
  assign _167_ = sc2mac_wt_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3608" *) sc2mac_wt_data43 : in_rt_wt_data_d1[351:344];
  assign _166_ = sc2mac_wt_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3598" *) sc2mac_wt_data42 : in_rt_wt_data_d1[343:336];
  assign _165_ = sc2mac_wt_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3588" *) sc2mac_wt_data41 : in_rt_wt_data_d1[335:328];
  assign _164_ = sc2mac_wt_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3578" *) sc2mac_wt_data40 : in_rt_wt_data_d1[327:320];
  assign _162_ = sc2mac_wt_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3568" *) sc2mac_wt_data39 : in_rt_wt_data_d1[319:312];
  assign _161_ = sc2mac_wt_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3558" *) sc2mac_wt_data38 : in_rt_wt_data_d1[311:304];
  assign _160_ = sc2mac_wt_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3548" *) sc2mac_wt_data37 : in_rt_wt_data_d1[303:296];
  assign _159_ = sc2mac_wt_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3538" *) sc2mac_wt_data36 : in_rt_wt_data_d1[295:288];
  assign _158_ = sc2mac_wt_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3528" *) sc2mac_wt_data35 : in_rt_wt_data_d1[287:280];
  assign _157_ = sc2mac_wt_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3518" *) sc2mac_wt_data34 : in_rt_wt_data_d1[279:272];
  assign _156_ = sc2mac_wt_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3508" *) sc2mac_wt_data33 : in_rt_wt_data_d1[271:264];
  assign _155_ = sc2mac_wt_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3498" *) sc2mac_wt_data32 : in_rt_wt_data_d1[263:256];
  assign _154_ = sc2mac_wt_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3488" *) sc2mac_wt_data31 : in_rt_wt_data_d1[255:248];
  assign _153_ = sc2mac_wt_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3478" *) sc2mac_wt_data30 : in_rt_wt_data_d1[247:240];
  assign _151_ = sc2mac_wt_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3468" *) sc2mac_wt_data29 : in_rt_wt_data_d1[239:232];
  assign _150_ = sc2mac_wt_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3458" *) sc2mac_wt_data28 : in_rt_wt_data_d1[231:224];
  assign _149_ = sc2mac_wt_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3448" *) sc2mac_wt_data27 : in_rt_wt_data_d1[223:216];
  assign _148_ = sc2mac_wt_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3438" *) sc2mac_wt_data26 : in_rt_wt_data_d1[215:208];
  assign _147_ = sc2mac_wt_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3428" *) sc2mac_wt_data25 : in_rt_wt_data_d1[207:200];
  assign _146_ = sc2mac_wt_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3418" *) sc2mac_wt_data24 : in_rt_wt_data_d1[199:192];
  assign _145_ = sc2mac_wt_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3408" *) sc2mac_wt_data23 : in_rt_wt_data_d1[191:184];
  assign _144_ = sc2mac_wt_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3398" *) sc2mac_wt_data22 : in_rt_wt_data_d1[183:176];
  assign _143_ = sc2mac_wt_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3388" *) sc2mac_wt_data21 : in_rt_wt_data_d1[175:168];
  assign _142_ = sc2mac_wt_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3378" *) sc2mac_wt_data20 : in_rt_wt_data_d1[167:160];
  assign _140_ = sc2mac_wt_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3368" *) sc2mac_wt_data19 : in_rt_wt_data_d1[159:152];
  assign _139_ = sc2mac_wt_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3358" *) sc2mac_wt_data18 : in_rt_wt_data_d1[151:144];
  assign _138_ = sc2mac_wt_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3348" *) sc2mac_wt_data17 : in_rt_wt_data_d1[143:136];
  assign _137_ = sc2mac_wt_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3338" *) sc2mac_wt_data16 : in_rt_wt_data_d1[135:128];
  assign _136_ = sc2mac_wt_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3328" *) sc2mac_wt_data15 : in_rt_wt_data_d1[127:120];
  assign _135_ = sc2mac_wt_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3318" *) sc2mac_wt_data14 : in_rt_wt_data_d1[119:112];
  assign _134_ = sc2mac_wt_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3308" *) sc2mac_wt_data13 : in_rt_wt_data_d1[111:104];
  assign _133_ = sc2mac_wt_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3298" *) sc2mac_wt_data12 : in_rt_wt_data_d1[103:96];
  assign _252_ = sc2mac_wt_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3288" *) sc2mac_wt_data11 : in_rt_wt_data_d1[95:88];
  assign _241_ = sc2mac_wt_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3278" *) sc2mac_wt_data10 : in_rt_wt_data_d1[87:80];
  assign _229_ = sc2mac_wt_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3268" *) sc2mac_wt_data9 : in_rt_wt_data_d1[79:72];
  assign _218_ = sc2mac_wt_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3258" *) sc2mac_wt_data8 : in_rt_wt_data_d1[71:64];
  assign _207_ = sc2mac_wt_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3248" *) sc2mac_wt_data7 : in_rt_wt_data_d1[63:56];
  assign _196_ = sc2mac_wt_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3238" *) sc2mac_wt_data6 : in_rt_wt_data_d1[55:48];
  assign _185_ = sc2mac_wt_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3228" *) sc2mac_wt_data5 : in_rt_wt_data_d1[47:40];
  assign _174_ = sc2mac_wt_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3218" *) sc2mac_wt_data4 : in_rt_wt_data_d1[39:32];
  assign _163_ = sc2mac_wt_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3208" *) sc2mac_wt_data3 : in_rt_wt_data_d1[31:24];
  assign _152_ = sc2mac_wt_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3198" *) sc2mac_wt_data2 : in_rt_wt_data_d1[23:16];
  assign _141_ = sc2mac_wt_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3188" *) sc2mac_wt_data1 : in_rt_wt_data_d1[15:8];
  assign _230_ = sc2mac_wt_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3178" *) sc2mac_wt_data0 : in_rt_wt_data_d1[7:0];
  assign _258_ = _261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3120" *) sc2mac_wt_mask : in_rt_wt_mask_d1;
  assign _259_ = _261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3059" *) sc2mac_wt_sel : in_rt_wt_sel_d1;
  assign _002_ = sc2mac_dat_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3039" *) sc2mac_dat_data127 : in_rt_dat_data_d1[1023:1016];
  assign _001_ = sc2mac_dat_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3029" *) sc2mac_dat_data126 : in_rt_dat_data_d1[1015:1008];
  assign _000_ = sc2mac_dat_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3019" *) sc2mac_dat_data125 : in_rt_dat_data_d1[1007:1000];
  assign _127_ = sc2mac_dat_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:3009" *) sc2mac_dat_data124 : in_rt_dat_data_d1[999:992];
  assign _126_ = sc2mac_dat_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2999" *) sc2mac_dat_data123 : in_rt_dat_data_d1[991:984];
  assign _125_ = sc2mac_dat_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2989" *) sc2mac_dat_data122 : in_rt_dat_data_d1[983:976];
  assign _124_ = sc2mac_dat_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2979" *) sc2mac_dat_data121 : in_rt_dat_data_d1[975:968];
  assign _123_ = sc2mac_dat_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2969" *) sc2mac_dat_data120 : in_rt_dat_data_d1[967:960];
  assign _121_ = sc2mac_dat_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2959" *) sc2mac_dat_data119 : in_rt_dat_data_d1[959:952];
  assign _120_ = sc2mac_dat_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2949" *) sc2mac_dat_data118 : in_rt_dat_data_d1[951:944];
  assign _119_ = sc2mac_dat_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2939" *) sc2mac_dat_data117 : in_rt_dat_data_d1[943:936];
  assign _118_ = sc2mac_dat_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2929" *) sc2mac_dat_data116 : in_rt_dat_data_d1[935:928];
  assign _117_ = sc2mac_dat_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2919" *) sc2mac_dat_data115 : in_rt_dat_data_d1[927:920];
  assign _116_ = sc2mac_dat_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2909" *) sc2mac_dat_data114 : in_rt_dat_data_d1[919:912];
  assign _115_ = sc2mac_dat_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2899" *) sc2mac_dat_data113 : in_rt_dat_data_d1[911:904];
  assign _114_ = sc2mac_dat_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2889" *) sc2mac_dat_data112 : in_rt_dat_data_d1[903:896];
  assign _113_ = sc2mac_dat_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2879" *) sc2mac_dat_data111 : in_rt_dat_data_d1[895:888];
  assign _112_ = sc2mac_dat_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2869" *) sc2mac_dat_data110 : in_rt_dat_data_d1[887:880];
  assign _110_ = sc2mac_dat_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2859" *) sc2mac_dat_data109 : in_rt_dat_data_d1[879:872];
  assign _109_ = sc2mac_dat_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2849" *) sc2mac_dat_data108 : in_rt_dat_data_d1[871:864];
  assign _108_ = sc2mac_dat_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2839" *) sc2mac_dat_data107 : in_rt_dat_data_d1[863:856];
  assign _107_ = sc2mac_dat_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2829" *) sc2mac_dat_data106 : in_rt_dat_data_d1[855:848];
  assign _106_ = sc2mac_dat_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2819" *) sc2mac_dat_data105 : in_rt_dat_data_d1[847:840];
  assign _105_ = sc2mac_dat_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2809" *) sc2mac_dat_data104 : in_rt_dat_data_d1[839:832];
  assign _104_ = sc2mac_dat_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2799" *) sc2mac_dat_data103 : in_rt_dat_data_d1[831:824];
  assign _103_ = sc2mac_dat_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2789" *) sc2mac_dat_data102 : in_rt_dat_data_d1[823:816];
  assign _102_ = sc2mac_dat_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2779" *) sc2mac_dat_data101 : in_rt_dat_data_d1[815:808];
  assign _101_ = sc2mac_dat_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2769" *) sc2mac_dat_data100 : in_rt_dat_data_d1[807:800];
  assign _098_ = sc2mac_dat_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2759" *) sc2mac_dat_data99 : in_rt_dat_data_d1[799:792];
  assign _097_ = sc2mac_dat_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2749" *) sc2mac_dat_data98 : in_rt_dat_data_d1[791:784];
  assign _096_ = sc2mac_dat_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2739" *) sc2mac_dat_data97 : in_rt_dat_data_d1[783:776];
  assign _095_ = sc2mac_dat_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2729" *) sc2mac_dat_data96 : in_rt_dat_data_d1[775:768];
  assign _094_ = sc2mac_dat_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2719" *) sc2mac_dat_data95 : in_rt_dat_data_d1[767:760];
  assign _093_ = sc2mac_dat_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2709" *) sc2mac_dat_data94 : in_rt_dat_data_d1[759:752];
  assign _092_ = sc2mac_dat_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2699" *) sc2mac_dat_data93 : in_rt_dat_data_d1[751:744];
  assign _091_ = sc2mac_dat_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2689" *) sc2mac_dat_data92 : in_rt_dat_data_d1[743:736];
  assign _090_ = sc2mac_dat_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2679" *) sc2mac_dat_data91 : in_rt_dat_data_d1[735:728];
  assign _089_ = sc2mac_dat_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2669" *) sc2mac_dat_data90 : in_rt_dat_data_d1[727:720];
  assign _087_ = sc2mac_dat_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2659" *) sc2mac_dat_data89 : in_rt_dat_data_d1[719:712];
  assign _086_ = sc2mac_dat_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2649" *) sc2mac_dat_data88 : in_rt_dat_data_d1[711:704];
  assign _085_ = sc2mac_dat_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2639" *) sc2mac_dat_data87 : in_rt_dat_data_d1[703:696];
  assign _084_ = sc2mac_dat_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2629" *) sc2mac_dat_data86 : in_rt_dat_data_d1[695:688];
  assign _083_ = sc2mac_dat_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2619" *) sc2mac_dat_data85 : in_rt_dat_data_d1[687:680];
  assign _082_ = sc2mac_dat_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2609" *) sc2mac_dat_data84 : in_rt_dat_data_d1[679:672];
  assign _081_ = sc2mac_dat_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2599" *) sc2mac_dat_data83 : in_rt_dat_data_d1[671:664];
  assign _080_ = sc2mac_dat_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2589" *) sc2mac_dat_data82 : in_rt_dat_data_d1[663:656];
  assign _079_ = sc2mac_dat_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2579" *) sc2mac_dat_data81 : in_rt_dat_data_d1[655:648];
  assign _078_ = sc2mac_dat_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2569" *) sc2mac_dat_data80 : in_rt_dat_data_d1[647:640];
  assign _076_ = sc2mac_dat_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2559" *) sc2mac_dat_data79 : in_rt_dat_data_d1[639:632];
  assign _075_ = sc2mac_dat_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2549" *) sc2mac_dat_data78 : in_rt_dat_data_d1[631:624];
  assign _074_ = sc2mac_dat_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2539" *) sc2mac_dat_data77 : in_rt_dat_data_d1[623:616];
  assign _073_ = sc2mac_dat_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2529" *) sc2mac_dat_data76 : in_rt_dat_data_d1[615:608];
  assign _072_ = sc2mac_dat_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2519" *) sc2mac_dat_data75 : in_rt_dat_data_d1[607:600];
  assign _071_ = sc2mac_dat_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2509" *) sc2mac_dat_data74 : in_rt_dat_data_d1[599:592];
  assign _070_ = sc2mac_dat_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2499" *) sc2mac_dat_data73 : in_rt_dat_data_d1[591:584];
  assign _069_ = sc2mac_dat_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2489" *) sc2mac_dat_data72 : in_rt_dat_data_d1[583:576];
  assign _068_ = sc2mac_dat_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2479" *) sc2mac_dat_data71 : in_rt_dat_data_d1[575:568];
  assign _067_ = sc2mac_dat_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2469" *) sc2mac_dat_data70 : in_rt_dat_data_d1[567:560];
  assign _065_ = sc2mac_dat_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2459" *) sc2mac_dat_data69 : in_rt_dat_data_d1[559:552];
  assign _064_ = sc2mac_dat_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2449" *) sc2mac_dat_data68 : in_rt_dat_data_d1[551:544];
  assign _063_ = sc2mac_dat_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2439" *) sc2mac_dat_data67 : in_rt_dat_data_d1[543:536];
  assign _062_ = sc2mac_dat_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2429" *) sc2mac_dat_data66 : in_rt_dat_data_d1[535:528];
  assign _061_ = sc2mac_dat_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2419" *) sc2mac_dat_data65 : in_rt_dat_data_d1[527:520];
  assign _060_ = sc2mac_dat_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2409" *) sc2mac_dat_data64 : in_rt_dat_data_d1[519:512];
  assign _059_ = sc2mac_dat_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2399" *) sc2mac_dat_data63 : in_rt_dat_data_d1[511:504];
  assign _058_ = sc2mac_dat_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2389" *) sc2mac_dat_data62 : in_rt_dat_data_d1[503:496];
  assign _057_ = sc2mac_dat_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2379" *) sc2mac_dat_data61 : in_rt_dat_data_d1[495:488];
  assign _056_ = sc2mac_dat_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2369" *) sc2mac_dat_data60 : in_rt_dat_data_d1[487:480];
  assign _054_ = sc2mac_dat_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2359" *) sc2mac_dat_data59 : in_rt_dat_data_d1[479:472];
  assign _053_ = sc2mac_dat_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2349" *) sc2mac_dat_data58 : in_rt_dat_data_d1[471:464];
  assign _052_ = sc2mac_dat_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2339" *) sc2mac_dat_data57 : in_rt_dat_data_d1[463:456];
  assign _051_ = sc2mac_dat_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2329" *) sc2mac_dat_data56 : in_rt_dat_data_d1[455:448];
  assign _050_ = sc2mac_dat_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2319" *) sc2mac_dat_data55 : in_rt_dat_data_d1[447:440];
  assign _049_ = sc2mac_dat_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2309" *) sc2mac_dat_data54 : in_rt_dat_data_d1[439:432];
  assign _048_ = sc2mac_dat_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2299" *) sc2mac_dat_data53 : in_rt_dat_data_d1[431:424];
  assign _047_ = sc2mac_dat_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2289" *) sc2mac_dat_data52 : in_rt_dat_data_d1[423:416];
  assign _046_ = sc2mac_dat_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2279" *) sc2mac_dat_data51 : in_rt_dat_data_d1[415:408];
  assign _045_ = sc2mac_dat_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2269" *) sc2mac_dat_data50 : in_rt_dat_data_d1[407:400];
  assign _043_ = sc2mac_dat_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2259" *) sc2mac_dat_data49 : in_rt_dat_data_d1[399:392];
  assign _042_ = sc2mac_dat_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2249" *) sc2mac_dat_data48 : in_rt_dat_data_d1[391:384];
  assign _041_ = sc2mac_dat_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2239" *) sc2mac_dat_data47 : in_rt_dat_data_d1[383:376];
  assign _040_ = sc2mac_dat_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2229" *) sc2mac_dat_data46 : in_rt_dat_data_d1[375:368];
  assign _039_ = sc2mac_dat_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2219" *) sc2mac_dat_data45 : in_rt_dat_data_d1[367:360];
  assign _038_ = sc2mac_dat_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2209" *) sc2mac_dat_data44 : in_rt_dat_data_d1[359:352];
  assign _037_ = sc2mac_dat_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2199" *) sc2mac_dat_data43 : in_rt_dat_data_d1[351:344];
  assign _036_ = sc2mac_dat_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2189" *) sc2mac_dat_data42 : in_rt_dat_data_d1[343:336];
  assign _035_ = sc2mac_dat_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2179" *) sc2mac_dat_data41 : in_rt_dat_data_d1[335:328];
  assign _034_ = sc2mac_dat_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2169" *) sc2mac_dat_data40 : in_rt_dat_data_d1[327:320];
  assign _032_ = sc2mac_dat_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2159" *) sc2mac_dat_data39 : in_rt_dat_data_d1[319:312];
  assign _031_ = sc2mac_dat_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2149" *) sc2mac_dat_data38 : in_rt_dat_data_d1[311:304];
  assign _030_ = sc2mac_dat_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2139" *) sc2mac_dat_data37 : in_rt_dat_data_d1[303:296];
  assign _029_ = sc2mac_dat_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2129" *) sc2mac_dat_data36 : in_rt_dat_data_d1[295:288];
  assign _028_ = sc2mac_dat_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2119" *) sc2mac_dat_data35 : in_rt_dat_data_d1[287:280];
  assign _027_ = sc2mac_dat_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2109" *) sc2mac_dat_data34 : in_rt_dat_data_d1[279:272];
  assign _026_ = sc2mac_dat_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2099" *) sc2mac_dat_data33 : in_rt_dat_data_d1[271:264];
  assign _025_ = sc2mac_dat_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2089" *) sc2mac_dat_data32 : in_rt_dat_data_d1[263:256];
  assign _024_ = sc2mac_dat_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2079" *) sc2mac_dat_data31 : in_rt_dat_data_d1[255:248];
  assign _023_ = sc2mac_dat_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2069" *) sc2mac_dat_data30 : in_rt_dat_data_d1[247:240];
  assign _021_ = sc2mac_dat_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2059" *) sc2mac_dat_data29 : in_rt_dat_data_d1[239:232];
  assign _020_ = sc2mac_dat_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2049" *) sc2mac_dat_data28 : in_rt_dat_data_d1[231:224];
  assign _019_ = sc2mac_dat_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2039" *) sc2mac_dat_data27 : in_rt_dat_data_d1[223:216];
  assign _018_ = sc2mac_dat_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2029" *) sc2mac_dat_data26 : in_rt_dat_data_d1[215:208];
  assign _017_ = sc2mac_dat_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2019" *) sc2mac_dat_data25 : in_rt_dat_data_d1[207:200];
  assign _016_ = sc2mac_dat_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:2009" *) sc2mac_dat_data24 : in_rt_dat_data_d1[199:192];
  assign _015_ = sc2mac_dat_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1999" *) sc2mac_dat_data23 : in_rt_dat_data_d1[191:184];
  assign _014_ = sc2mac_dat_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1989" *) sc2mac_dat_data22 : in_rt_dat_data_d1[183:176];
  assign _013_ = sc2mac_dat_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1979" *) sc2mac_dat_data21 : in_rt_dat_data_d1[175:168];
  assign _012_ = sc2mac_dat_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1969" *) sc2mac_dat_data20 : in_rt_dat_data_d1[167:160];
  assign _010_ = sc2mac_dat_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1959" *) sc2mac_dat_data19 : in_rt_dat_data_d1[159:152];
  assign _009_ = sc2mac_dat_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1949" *) sc2mac_dat_data18 : in_rt_dat_data_d1[151:144];
  assign _008_ = sc2mac_dat_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1939" *) sc2mac_dat_data17 : in_rt_dat_data_d1[143:136];
  assign _007_ = sc2mac_dat_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1929" *) sc2mac_dat_data16 : in_rt_dat_data_d1[135:128];
  assign _006_ = sc2mac_dat_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1919" *) sc2mac_dat_data15 : in_rt_dat_data_d1[127:120];
  assign _005_ = sc2mac_dat_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1909" *) sc2mac_dat_data14 : in_rt_dat_data_d1[119:112];
  assign _004_ = sc2mac_dat_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1899" *) sc2mac_dat_data13 : in_rt_dat_data_d1[111:104];
  assign _003_ = sc2mac_dat_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1889" *) sc2mac_dat_data12 : in_rt_dat_data_d1[103:96];
  assign _122_ = sc2mac_dat_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1879" *) sc2mac_dat_data11 : in_rt_dat_data_d1[95:88];
  assign _111_ = sc2mac_dat_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1869" *) sc2mac_dat_data10 : in_rt_dat_data_d1[87:80];
  assign _099_ = sc2mac_dat_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1859" *) sc2mac_dat_data9 : in_rt_dat_data_d1[79:72];
  assign _088_ = sc2mac_dat_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1849" *) sc2mac_dat_data8 : in_rt_dat_data_d1[71:64];
  assign _077_ = sc2mac_dat_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1839" *) sc2mac_dat_data7 : in_rt_dat_data_d1[63:56];
  assign _066_ = sc2mac_dat_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1829" *) sc2mac_dat_data6 : in_rt_dat_data_d1[55:48];
  assign _055_ = sc2mac_dat_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1819" *) sc2mac_dat_data5 : in_rt_dat_data_d1[47:40];
  assign _044_ = sc2mac_dat_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1809" *) sc2mac_dat_data4 : in_rt_dat_data_d1[39:32];
  assign _033_ = sc2mac_dat_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1799" *) sc2mac_dat_data3 : in_rt_dat_data_d1[31:24];
  assign _022_ = sc2mac_dat_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1789" *) sc2mac_dat_data2 : in_rt_dat_data_d1[23:16];
  assign _011_ = sc2mac_dat_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1779" *) sc2mac_dat_data1 : in_rt_dat_data_d1[15:8];
  assign _100_ = sc2mac_dat_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1769" *) sc2mac_dat_data0 : in_rt_dat_data_d1[7:0];
  assign _129_ = _260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1711" *) sc2mac_dat_pd : in_rt_dat_pd_d1;
  assign _128_ = _260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_rt_in.v:1650" *) sc2mac_dat_mask : in_rt_dat_mask_d1;
  assign in_dat_data = in_rt_dat_data_d1;
  assign in_dat_data0 = in_rt_dat_data_d1[7:0];
  assign in_dat_data1 = in_rt_dat_data_d1[15:8];
  assign in_dat_data10 = in_rt_dat_data_d1[87:80];
  assign in_dat_data100 = in_rt_dat_data_d1[807:800];
  assign in_dat_data101 = in_rt_dat_data_d1[815:808];
  assign in_dat_data102 = in_rt_dat_data_d1[823:816];
  assign in_dat_data103 = in_rt_dat_data_d1[831:824];
  assign in_dat_data104 = in_rt_dat_data_d1[839:832];
  assign in_dat_data105 = in_rt_dat_data_d1[847:840];
  assign in_dat_data106 = in_rt_dat_data_d1[855:848];
  assign in_dat_data107 = in_rt_dat_data_d1[863:856];
  assign in_dat_data108 = in_rt_dat_data_d1[871:864];
  assign in_dat_data109 = in_rt_dat_data_d1[879:872];
  assign in_dat_data11 = in_rt_dat_data_d1[95:88];
  assign in_dat_data110 = in_rt_dat_data_d1[887:880];
  assign in_dat_data111 = in_rt_dat_data_d1[895:888];
  assign in_dat_data112 = in_rt_dat_data_d1[903:896];
  assign in_dat_data113 = in_rt_dat_data_d1[911:904];
  assign in_dat_data114 = in_rt_dat_data_d1[919:912];
  assign in_dat_data115 = in_rt_dat_data_d1[927:920];
  assign in_dat_data116 = in_rt_dat_data_d1[935:928];
  assign in_dat_data117 = in_rt_dat_data_d1[943:936];
  assign in_dat_data118 = in_rt_dat_data_d1[951:944];
  assign in_dat_data119 = in_rt_dat_data_d1[959:952];
  assign in_dat_data12 = in_rt_dat_data_d1[103:96];
  assign in_dat_data120 = in_rt_dat_data_d1[967:960];
  assign in_dat_data121 = in_rt_dat_data_d1[975:968];
  assign in_dat_data122 = in_rt_dat_data_d1[983:976];
  assign in_dat_data123 = in_rt_dat_data_d1[991:984];
  assign in_dat_data124 = in_rt_dat_data_d1[999:992];
  assign in_dat_data125 = in_rt_dat_data_d1[1007:1000];
  assign in_dat_data126 = in_rt_dat_data_d1[1015:1008];
  assign in_dat_data127 = in_rt_dat_data_d1[1023:1016];
  assign in_dat_data13 = in_rt_dat_data_d1[111:104];
  assign in_dat_data14 = in_rt_dat_data_d1[119:112];
  assign in_dat_data15 = in_rt_dat_data_d1[127:120];
  assign in_dat_data16 = in_rt_dat_data_d1[135:128];
  assign in_dat_data17 = in_rt_dat_data_d1[143:136];
  assign in_dat_data18 = in_rt_dat_data_d1[151:144];
  assign in_dat_data19 = in_rt_dat_data_d1[159:152];
  assign in_dat_data2 = in_rt_dat_data_d1[23:16];
  assign in_dat_data20 = in_rt_dat_data_d1[167:160];
  assign in_dat_data21 = in_rt_dat_data_d1[175:168];
  assign in_dat_data22 = in_rt_dat_data_d1[183:176];
  assign in_dat_data23 = in_rt_dat_data_d1[191:184];
  assign in_dat_data24 = in_rt_dat_data_d1[199:192];
  assign in_dat_data25 = in_rt_dat_data_d1[207:200];
  assign in_dat_data26 = in_rt_dat_data_d1[215:208];
  assign in_dat_data27 = in_rt_dat_data_d1[223:216];
  assign in_dat_data28 = in_rt_dat_data_d1[231:224];
  assign in_dat_data29 = in_rt_dat_data_d1[239:232];
  assign in_dat_data3 = in_rt_dat_data_d1[31:24];
  assign in_dat_data30 = in_rt_dat_data_d1[247:240];
  assign in_dat_data31 = in_rt_dat_data_d1[255:248];
  assign in_dat_data32 = in_rt_dat_data_d1[263:256];
  assign in_dat_data33 = in_rt_dat_data_d1[271:264];
  assign in_dat_data34 = in_rt_dat_data_d1[279:272];
  assign in_dat_data35 = in_rt_dat_data_d1[287:280];
  assign in_dat_data36 = in_rt_dat_data_d1[295:288];
  assign in_dat_data37 = in_rt_dat_data_d1[303:296];
  assign in_dat_data38 = in_rt_dat_data_d1[311:304];
  assign in_dat_data39 = in_rt_dat_data_d1[319:312];
  assign in_dat_data4 = in_rt_dat_data_d1[39:32];
  assign in_dat_data40 = in_rt_dat_data_d1[327:320];
  assign in_dat_data41 = in_rt_dat_data_d1[335:328];
  assign in_dat_data42 = in_rt_dat_data_d1[343:336];
  assign in_dat_data43 = in_rt_dat_data_d1[351:344];
  assign in_dat_data44 = in_rt_dat_data_d1[359:352];
  assign in_dat_data45 = in_rt_dat_data_d1[367:360];
  assign in_dat_data46 = in_rt_dat_data_d1[375:368];
  assign in_dat_data47 = in_rt_dat_data_d1[383:376];
  assign in_dat_data48 = in_rt_dat_data_d1[391:384];
  assign in_dat_data49 = in_rt_dat_data_d1[399:392];
  assign in_dat_data5 = in_rt_dat_data_d1[47:40];
  assign in_dat_data50 = in_rt_dat_data_d1[407:400];
  assign in_dat_data51 = in_rt_dat_data_d1[415:408];
  assign in_dat_data52 = in_rt_dat_data_d1[423:416];
  assign in_dat_data53 = in_rt_dat_data_d1[431:424];
  assign in_dat_data54 = in_rt_dat_data_d1[439:432];
  assign in_dat_data55 = in_rt_dat_data_d1[447:440];
  assign in_dat_data56 = in_rt_dat_data_d1[455:448];
  assign in_dat_data57 = in_rt_dat_data_d1[463:456];
  assign in_dat_data58 = in_rt_dat_data_d1[471:464];
  assign in_dat_data59 = in_rt_dat_data_d1[479:472];
  assign in_dat_data6 = in_rt_dat_data_d1[55:48];
  assign in_dat_data60 = in_rt_dat_data_d1[487:480];
  assign in_dat_data61 = in_rt_dat_data_d1[495:488];
  assign in_dat_data62 = in_rt_dat_data_d1[503:496];
  assign in_dat_data63 = in_rt_dat_data_d1[511:504];
  assign in_dat_data64 = in_rt_dat_data_d1[519:512];
  assign in_dat_data65 = in_rt_dat_data_d1[527:520];
  assign in_dat_data66 = in_rt_dat_data_d1[535:528];
  assign in_dat_data67 = in_rt_dat_data_d1[543:536];
  assign in_dat_data68 = in_rt_dat_data_d1[551:544];
  assign in_dat_data69 = in_rt_dat_data_d1[559:552];
  assign in_dat_data7 = in_rt_dat_data_d1[63:56];
  assign in_dat_data70 = in_rt_dat_data_d1[567:560];
  assign in_dat_data71 = in_rt_dat_data_d1[575:568];
  assign in_dat_data72 = in_rt_dat_data_d1[583:576];
  assign in_dat_data73 = in_rt_dat_data_d1[591:584];
  assign in_dat_data74 = in_rt_dat_data_d1[599:592];
  assign in_dat_data75 = in_rt_dat_data_d1[607:600];
  assign in_dat_data76 = in_rt_dat_data_d1[615:608];
  assign in_dat_data77 = in_rt_dat_data_d1[623:616];
  assign in_dat_data78 = in_rt_dat_data_d1[631:624];
  assign in_dat_data79 = in_rt_dat_data_d1[639:632];
  assign in_dat_data8 = in_rt_dat_data_d1[71:64];
  assign in_dat_data80 = in_rt_dat_data_d1[647:640];
  assign in_dat_data81 = in_rt_dat_data_d1[655:648];
  assign in_dat_data82 = in_rt_dat_data_d1[663:656];
  assign in_dat_data83 = in_rt_dat_data_d1[671:664];
  assign in_dat_data84 = in_rt_dat_data_d1[679:672];
  assign in_dat_data85 = in_rt_dat_data_d1[687:680];
  assign in_dat_data86 = in_rt_dat_data_d1[695:688];
  assign in_dat_data87 = in_rt_dat_data_d1[703:696];
  assign in_dat_data88 = in_rt_dat_data_d1[711:704];
  assign in_dat_data89 = in_rt_dat_data_d1[719:712];
  assign in_dat_data9 = in_rt_dat_data_d1[79:72];
  assign in_dat_data90 = in_rt_dat_data_d1[727:720];
  assign in_dat_data91 = in_rt_dat_data_d1[735:728];
  assign in_dat_data92 = in_rt_dat_data_d1[743:736];
  assign in_dat_data93 = in_rt_dat_data_d1[751:744];
  assign in_dat_data94 = in_rt_dat_data_d1[759:752];
  assign in_dat_data95 = in_rt_dat_data_d1[767:760];
  assign in_dat_data96 = in_rt_dat_data_d1[775:768];
  assign in_dat_data97 = in_rt_dat_data_d1[783:776];
  assign in_dat_data98 = in_rt_dat_data_d1[791:784];
  assign in_dat_data99 = in_rt_dat_data_d1[799:792];
  assign in_dat_mask = in_rt_dat_mask_d1;
  assign in_dat_pd = in_rt_dat_pd_d1;
  assign in_dat_pvld = in_rt_dat_pvld_d1;
  assign in_dat_stripe_end = in_rt_dat_pd_d1[6];
  assign in_dat_stripe_st = in_rt_dat_pd_d1[5];
  assign in_rt_dat_data_d0 = { sc2mac_dat_data127, sc2mac_dat_data126, sc2mac_dat_data125, sc2mac_dat_data124, sc2mac_dat_data123, sc2mac_dat_data122, sc2mac_dat_data121, sc2mac_dat_data120, sc2mac_dat_data119, sc2mac_dat_data118, sc2mac_dat_data117, sc2mac_dat_data116, sc2mac_dat_data115, sc2mac_dat_data114, sc2mac_dat_data113, sc2mac_dat_data112, sc2mac_dat_data111, sc2mac_dat_data110, sc2mac_dat_data109, sc2mac_dat_data108, sc2mac_dat_data107, sc2mac_dat_data106, sc2mac_dat_data105, sc2mac_dat_data104, sc2mac_dat_data103, sc2mac_dat_data102, sc2mac_dat_data101, sc2mac_dat_data100, sc2mac_dat_data99, sc2mac_dat_data98, sc2mac_dat_data97, sc2mac_dat_data96, sc2mac_dat_data95, sc2mac_dat_data94, sc2mac_dat_data93, sc2mac_dat_data92, sc2mac_dat_data91, sc2mac_dat_data90, sc2mac_dat_data89, sc2mac_dat_data88, sc2mac_dat_data87, sc2mac_dat_data86, sc2mac_dat_data85, sc2mac_dat_data84, sc2mac_dat_data83, sc2mac_dat_data82, sc2mac_dat_data81, sc2mac_dat_data80, sc2mac_dat_data79, sc2mac_dat_data78, sc2mac_dat_data77, sc2mac_dat_data76, sc2mac_dat_data75, sc2mac_dat_data74, sc2mac_dat_data73, sc2mac_dat_data72, sc2mac_dat_data71, sc2mac_dat_data70, sc2mac_dat_data69, sc2mac_dat_data68, sc2mac_dat_data67, sc2mac_dat_data66, sc2mac_dat_data65, sc2mac_dat_data64, sc2mac_dat_data63, sc2mac_dat_data62, sc2mac_dat_data61, sc2mac_dat_data60, sc2mac_dat_data59, sc2mac_dat_data58, sc2mac_dat_data57, sc2mac_dat_data56, sc2mac_dat_data55, sc2mac_dat_data54, sc2mac_dat_data53, sc2mac_dat_data52, sc2mac_dat_data51, sc2mac_dat_data50, sc2mac_dat_data49, sc2mac_dat_data48, sc2mac_dat_data47, sc2mac_dat_data46, sc2mac_dat_data45, sc2mac_dat_data44, sc2mac_dat_data43, sc2mac_dat_data42, sc2mac_dat_data41, sc2mac_dat_data40, sc2mac_dat_data39, sc2mac_dat_data38, sc2mac_dat_data37, sc2mac_dat_data36, sc2mac_dat_data35, sc2mac_dat_data34, sc2mac_dat_data33, sc2mac_dat_data32, sc2mac_dat_data31, sc2mac_dat_data30, sc2mac_dat_data29, sc2mac_dat_data28, sc2mac_dat_data27, sc2mac_dat_data26, sc2mac_dat_data25, sc2mac_dat_data24, sc2mac_dat_data23, sc2mac_dat_data22, sc2mac_dat_data21, sc2mac_dat_data20, sc2mac_dat_data19, sc2mac_dat_data18, sc2mac_dat_data17, sc2mac_dat_data16, sc2mac_dat_data15, sc2mac_dat_data14, sc2mac_dat_data13, sc2mac_dat_data12, sc2mac_dat_data11, sc2mac_dat_data10, sc2mac_dat_data9, sc2mac_dat_data8, sc2mac_dat_data7, sc2mac_dat_data6, sc2mac_dat_data5, sc2mac_dat_data4, sc2mac_dat_data3, sc2mac_dat_data2, sc2mac_dat_data1, sc2mac_dat_data0 };
  assign in_rt_dat_mask_d0 = sc2mac_dat_mask;
  assign in_rt_dat_pd_d0 = sc2mac_dat_pd;
  assign in_rt_dat_pvld_d0 = sc2mac_dat_pvld;
  assign in_rt_wt_data_d0 = { sc2mac_wt_data127, sc2mac_wt_data126, sc2mac_wt_data125, sc2mac_wt_data124, sc2mac_wt_data123, sc2mac_wt_data122, sc2mac_wt_data121, sc2mac_wt_data120, sc2mac_wt_data119, sc2mac_wt_data118, sc2mac_wt_data117, sc2mac_wt_data116, sc2mac_wt_data115, sc2mac_wt_data114, sc2mac_wt_data113, sc2mac_wt_data112, sc2mac_wt_data111, sc2mac_wt_data110, sc2mac_wt_data109, sc2mac_wt_data108, sc2mac_wt_data107, sc2mac_wt_data106, sc2mac_wt_data105, sc2mac_wt_data104, sc2mac_wt_data103, sc2mac_wt_data102, sc2mac_wt_data101, sc2mac_wt_data100, sc2mac_wt_data99, sc2mac_wt_data98, sc2mac_wt_data97, sc2mac_wt_data96, sc2mac_wt_data95, sc2mac_wt_data94, sc2mac_wt_data93, sc2mac_wt_data92, sc2mac_wt_data91, sc2mac_wt_data90, sc2mac_wt_data89, sc2mac_wt_data88, sc2mac_wt_data87, sc2mac_wt_data86, sc2mac_wt_data85, sc2mac_wt_data84, sc2mac_wt_data83, sc2mac_wt_data82, sc2mac_wt_data81, sc2mac_wt_data80, sc2mac_wt_data79, sc2mac_wt_data78, sc2mac_wt_data77, sc2mac_wt_data76, sc2mac_wt_data75, sc2mac_wt_data74, sc2mac_wt_data73, sc2mac_wt_data72, sc2mac_wt_data71, sc2mac_wt_data70, sc2mac_wt_data69, sc2mac_wt_data68, sc2mac_wt_data67, sc2mac_wt_data66, sc2mac_wt_data65, sc2mac_wt_data64, sc2mac_wt_data63, sc2mac_wt_data62, sc2mac_wt_data61, sc2mac_wt_data60, sc2mac_wt_data59, sc2mac_wt_data58, sc2mac_wt_data57, sc2mac_wt_data56, sc2mac_wt_data55, sc2mac_wt_data54, sc2mac_wt_data53, sc2mac_wt_data52, sc2mac_wt_data51, sc2mac_wt_data50, sc2mac_wt_data49, sc2mac_wt_data48, sc2mac_wt_data47, sc2mac_wt_data46, sc2mac_wt_data45, sc2mac_wt_data44, sc2mac_wt_data43, sc2mac_wt_data42, sc2mac_wt_data41, sc2mac_wt_data40, sc2mac_wt_data39, sc2mac_wt_data38, sc2mac_wt_data37, sc2mac_wt_data36, sc2mac_wt_data35, sc2mac_wt_data34, sc2mac_wt_data33, sc2mac_wt_data32, sc2mac_wt_data31, sc2mac_wt_data30, sc2mac_wt_data29, sc2mac_wt_data28, sc2mac_wt_data27, sc2mac_wt_data26, sc2mac_wt_data25, sc2mac_wt_data24, sc2mac_wt_data23, sc2mac_wt_data22, sc2mac_wt_data21, sc2mac_wt_data20, sc2mac_wt_data19, sc2mac_wt_data18, sc2mac_wt_data17, sc2mac_wt_data16, sc2mac_wt_data15, sc2mac_wt_data14, sc2mac_wt_data13, sc2mac_wt_data12, sc2mac_wt_data11, sc2mac_wt_data10, sc2mac_wt_data9, sc2mac_wt_data8, sc2mac_wt_data7, sc2mac_wt_data6, sc2mac_wt_data5, sc2mac_wt_data4, sc2mac_wt_data3, sc2mac_wt_data2, sc2mac_wt_data1, sc2mac_wt_data0 };
  assign in_rt_wt_mask_d0 = sc2mac_wt_mask;
  assign in_rt_wt_pvld_d0 = sc2mac_wt_pvld;
  assign in_rt_wt_sel_d0 = sc2mac_wt_sel;
  assign in_wt_data = in_rt_wt_data_d1;
  assign in_wt_data0 = in_rt_wt_data_d1[7:0];
  assign in_wt_data1 = in_rt_wt_data_d1[15:8];
  assign in_wt_data10 = in_rt_wt_data_d1[87:80];
  assign in_wt_data100 = in_rt_wt_data_d1[807:800];
  assign in_wt_data101 = in_rt_wt_data_d1[815:808];
  assign in_wt_data102 = in_rt_wt_data_d1[823:816];
  assign in_wt_data103 = in_rt_wt_data_d1[831:824];
  assign in_wt_data104 = in_rt_wt_data_d1[839:832];
  assign in_wt_data105 = in_rt_wt_data_d1[847:840];
  assign in_wt_data106 = in_rt_wt_data_d1[855:848];
  assign in_wt_data107 = in_rt_wt_data_d1[863:856];
  assign in_wt_data108 = in_rt_wt_data_d1[871:864];
  assign in_wt_data109 = in_rt_wt_data_d1[879:872];
  assign in_wt_data11 = in_rt_wt_data_d1[95:88];
  assign in_wt_data110 = in_rt_wt_data_d1[887:880];
  assign in_wt_data111 = in_rt_wt_data_d1[895:888];
  assign in_wt_data112 = in_rt_wt_data_d1[903:896];
  assign in_wt_data113 = in_rt_wt_data_d1[911:904];
  assign in_wt_data114 = in_rt_wt_data_d1[919:912];
  assign in_wt_data115 = in_rt_wt_data_d1[927:920];
  assign in_wt_data116 = in_rt_wt_data_d1[935:928];
  assign in_wt_data117 = in_rt_wt_data_d1[943:936];
  assign in_wt_data118 = in_rt_wt_data_d1[951:944];
  assign in_wt_data119 = in_rt_wt_data_d1[959:952];
  assign in_wt_data12 = in_rt_wt_data_d1[103:96];
  assign in_wt_data120 = in_rt_wt_data_d1[967:960];
  assign in_wt_data121 = in_rt_wt_data_d1[975:968];
  assign in_wt_data122 = in_rt_wt_data_d1[983:976];
  assign in_wt_data123 = in_rt_wt_data_d1[991:984];
  assign in_wt_data124 = in_rt_wt_data_d1[999:992];
  assign in_wt_data125 = in_rt_wt_data_d1[1007:1000];
  assign in_wt_data126 = in_rt_wt_data_d1[1015:1008];
  assign in_wt_data127 = in_rt_wt_data_d1[1023:1016];
  assign in_wt_data13 = in_rt_wt_data_d1[111:104];
  assign in_wt_data14 = in_rt_wt_data_d1[119:112];
  assign in_wt_data15 = in_rt_wt_data_d1[127:120];
  assign in_wt_data16 = in_rt_wt_data_d1[135:128];
  assign in_wt_data17 = in_rt_wt_data_d1[143:136];
  assign in_wt_data18 = in_rt_wt_data_d1[151:144];
  assign in_wt_data19 = in_rt_wt_data_d1[159:152];
  assign in_wt_data2 = in_rt_wt_data_d1[23:16];
  assign in_wt_data20 = in_rt_wt_data_d1[167:160];
  assign in_wt_data21 = in_rt_wt_data_d1[175:168];
  assign in_wt_data22 = in_rt_wt_data_d1[183:176];
  assign in_wt_data23 = in_rt_wt_data_d1[191:184];
  assign in_wt_data24 = in_rt_wt_data_d1[199:192];
  assign in_wt_data25 = in_rt_wt_data_d1[207:200];
  assign in_wt_data26 = in_rt_wt_data_d1[215:208];
  assign in_wt_data27 = in_rt_wt_data_d1[223:216];
  assign in_wt_data28 = in_rt_wt_data_d1[231:224];
  assign in_wt_data29 = in_rt_wt_data_d1[239:232];
  assign in_wt_data3 = in_rt_wt_data_d1[31:24];
  assign in_wt_data30 = in_rt_wt_data_d1[247:240];
  assign in_wt_data31 = in_rt_wt_data_d1[255:248];
  assign in_wt_data32 = in_rt_wt_data_d1[263:256];
  assign in_wt_data33 = in_rt_wt_data_d1[271:264];
  assign in_wt_data34 = in_rt_wt_data_d1[279:272];
  assign in_wt_data35 = in_rt_wt_data_d1[287:280];
  assign in_wt_data36 = in_rt_wt_data_d1[295:288];
  assign in_wt_data37 = in_rt_wt_data_d1[303:296];
  assign in_wt_data38 = in_rt_wt_data_d1[311:304];
  assign in_wt_data39 = in_rt_wt_data_d1[319:312];
  assign in_wt_data4 = in_rt_wt_data_d1[39:32];
  assign in_wt_data40 = in_rt_wt_data_d1[327:320];
  assign in_wt_data41 = in_rt_wt_data_d1[335:328];
  assign in_wt_data42 = in_rt_wt_data_d1[343:336];
  assign in_wt_data43 = in_rt_wt_data_d1[351:344];
  assign in_wt_data44 = in_rt_wt_data_d1[359:352];
  assign in_wt_data45 = in_rt_wt_data_d1[367:360];
  assign in_wt_data46 = in_rt_wt_data_d1[375:368];
  assign in_wt_data47 = in_rt_wt_data_d1[383:376];
  assign in_wt_data48 = in_rt_wt_data_d1[391:384];
  assign in_wt_data49 = in_rt_wt_data_d1[399:392];
  assign in_wt_data5 = in_rt_wt_data_d1[47:40];
  assign in_wt_data50 = in_rt_wt_data_d1[407:400];
  assign in_wt_data51 = in_rt_wt_data_d1[415:408];
  assign in_wt_data52 = in_rt_wt_data_d1[423:416];
  assign in_wt_data53 = in_rt_wt_data_d1[431:424];
  assign in_wt_data54 = in_rt_wt_data_d1[439:432];
  assign in_wt_data55 = in_rt_wt_data_d1[447:440];
  assign in_wt_data56 = in_rt_wt_data_d1[455:448];
  assign in_wt_data57 = in_rt_wt_data_d1[463:456];
  assign in_wt_data58 = in_rt_wt_data_d1[471:464];
  assign in_wt_data59 = in_rt_wt_data_d1[479:472];
  assign in_wt_data6 = in_rt_wt_data_d1[55:48];
  assign in_wt_data60 = in_rt_wt_data_d1[487:480];
  assign in_wt_data61 = in_rt_wt_data_d1[495:488];
  assign in_wt_data62 = in_rt_wt_data_d1[503:496];
  assign in_wt_data63 = in_rt_wt_data_d1[511:504];
  assign in_wt_data64 = in_rt_wt_data_d1[519:512];
  assign in_wt_data65 = in_rt_wt_data_d1[527:520];
  assign in_wt_data66 = in_rt_wt_data_d1[535:528];
  assign in_wt_data67 = in_rt_wt_data_d1[543:536];
  assign in_wt_data68 = in_rt_wt_data_d1[551:544];
  assign in_wt_data69 = in_rt_wt_data_d1[559:552];
  assign in_wt_data7 = in_rt_wt_data_d1[63:56];
  assign in_wt_data70 = in_rt_wt_data_d1[567:560];
  assign in_wt_data71 = in_rt_wt_data_d1[575:568];
  assign in_wt_data72 = in_rt_wt_data_d1[583:576];
  assign in_wt_data73 = in_rt_wt_data_d1[591:584];
  assign in_wt_data74 = in_rt_wt_data_d1[599:592];
  assign in_wt_data75 = in_rt_wt_data_d1[607:600];
  assign in_wt_data76 = in_rt_wt_data_d1[615:608];
  assign in_wt_data77 = in_rt_wt_data_d1[623:616];
  assign in_wt_data78 = in_rt_wt_data_d1[631:624];
  assign in_wt_data79 = in_rt_wt_data_d1[639:632];
  assign in_wt_data8 = in_rt_wt_data_d1[71:64];
  assign in_wt_data80 = in_rt_wt_data_d1[647:640];
  assign in_wt_data81 = in_rt_wt_data_d1[655:648];
  assign in_wt_data82 = in_rt_wt_data_d1[663:656];
  assign in_wt_data83 = in_rt_wt_data_d1[671:664];
  assign in_wt_data84 = in_rt_wt_data_d1[679:672];
  assign in_wt_data85 = in_rt_wt_data_d1[687:680];
  assign in_wt_data86 = in_rt_wt_data_d1[695:688];
  assign in_wt_data87 = in_rt_wt_data_d1[703:696];
  assign in_wt_data88 = in_rt_wt_data_d1[711:704];
  assign in_wt_data89 = in_rt_wt_data_d1[719:712];
  assign in_wt_data9 = in_rt_wt_data_d1[79:72];
  assign in_wt_data90 = in_rt_wt_data_d1[727:720];
  assign in_wt_data91 = in_rt_wt_data_d1[735:728];
  assign in_wt_data92 = in_rt_wt_data_d1[743:736];
  assign in_wt_data93 = in_rt_wt_data_d1[751:744];
  assign in_wt_data94 = in_rt_wt_data_d1[759:752];
  assign in_wt_data95 = in_rt_wt_data_d1[767:760];
  assign in_wt_data96 = in_rt_wt_data_d1[775:768];
  assign in_wt_data97 = in_rt_wt_data_d1[783:776];
  assign in_wt_data98 = in_rt_wt_data_d1[791:784];
  assign in_wt_data99 = in_rt_wt_data_d1[799:792];
  assign in_wt_mask = in_rt_wt_mask_d1;
  assign in_wt_pvld = in_rt_wt_pvld_d1;
  assign in_wt_sel = in_rt_wt_sel_d1;
endmodule
