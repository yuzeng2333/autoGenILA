module NV_BLKBOX_SRC0_X(Y);
  (* src = "./vmod/vlibs/NV_BLKBOX_SRC0_X.v:12" *)
  output Y;
  assign Y = 1'b0;
endmodule
