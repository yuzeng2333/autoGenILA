module CDMA_chn_data_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:369" *)
  input in_0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:370" *)
  output outsig;
  assign outsig = in_0;
endmodule
