module UINT16_TO_FP17_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_uint16_to_fp17.v:201" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_uint16_to_fp17.v:202" *)
  output outsig;
  assign outsig = in_0;
endmodule
