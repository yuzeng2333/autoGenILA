module \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=8\width=1 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:78" *)
  output d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:79" *)
  input z;
  assign d = z;
endmodule
