module \$paramod\SDP_C_mgc_in_wire_v1\rscid=5\width=2 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:78" *)
  output [1:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:79" *)
  input [1:0] z;
  assign d = z;
endmodule
