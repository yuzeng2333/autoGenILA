module NV_NVDLA_CDMA_IMG_pack(nvdla_core_clk, nvdla_core_rstn, img2sbuf_p0_rd_data, img2sbuf_p1_rd_data, is_running, layer_st, pixel_bank, pixel_data_expand, pixel_data_shrink, pixel_early_end, pixel_packed_10b, pixel_planar, pixel_planar0_sft, pixel_planar1_sft, pixel_precision, pixel_uint, reg2dp_datain_channel, reg2dp_datain_width, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_pad_left, reg2dp_pad_right, sg2pack_data_entries, sg2pack_entry_end, sg2pack_entry_mid, sg2pack_entry_st, sg2pack_height_total, sg2pack_img_pd, sg2pack_img_pvld, sg2pack_mn_enable, sg2pack_sub_h_end, sg2pack_sub_h_mid, sg2pack_sub_h_st, status2dma_wr_idx, img2cvt_dat_wr_addr, img2cvt_dat_wr_data, img2cvt_dat_wr_en, img2cvt_dat_wr_hsel, img2cvt_dat_wr_info_pd, img2cvt_dat_wr_pad_mask, img2cvt_mn_wr_data, img2sbuf_p0_rd_addr, img2sbuf_p0_rd_en, img2sbuf_p1_rd_addr, img2sbuf_p1_rd_en, img2status_dat_entries, img2status_dat_slices, img2status_dat_updt, pack_is_done, sg2pack_img_prdy);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1125" *)
  wire [5:0] _0000_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2795" *)
  wire [13:0] _0001_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3039" *)
  wire [2:0] _0002_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1186" *)
  wire [5:0] _0003_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2856" *)
  wire [13:0] _0004_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3100" *)
  wire [2:0] _0005_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:637" *)
  wire [13:0] _0006_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:698" *)
  wire [13:0] _0007_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:759" *)
  wire [4:0] _0008_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:820" *)
  wire [4:0] _0009_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6479" *)
  wire [63:0] _0010_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7076" *)
  wire [63:0] _0011_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:576" *)
  wire [4:0] _0012_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7269" *)
  wire [511:0] _0013_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7259" *)
  wire [511:0] _0014_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7996" *)
  wire [11:0] _0015_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8278" *)
  wire [11:0] _0016_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6672" *)
  wire [511:0] _0017_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6662" *)
  wire [511:0] _0018_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8339" *)
  wire [3:0] _0019_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5880" *)
  wire _0020_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5819" *)
  wire _0021_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8057" *)
  wire _0022_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5636" *)
  wire [3:0] _0023_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5697" *)
  wire _0024_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6743" *)
  wire [63:0] _0025_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6682" *)
  wire [63:0] _0026_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5575" *)
  wire [2:0] _0027_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5758" *)
  wire _0028_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5349" *)
  wire _0029_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5410" *)
  wire _0030_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5227" *)
  wire _0031_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5288" *)
  wire _0032_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6296" *)
  wire [511:0] _0033_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5105" *)
  wire [2:0] _0034_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5166" *)
  wire _0035_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7344" *)
  wire [11:0] _0036_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5502" *)
  wire [1:0] _0037_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7517" *)
  wire [11:0] _0038_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7703" *)
  wire [13:0] _0039_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7764" *)
  wire [13:0] _0040_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3588" *)
  wire _0041_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4448" *)
  wire _0042_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4922" *)
  wire _0043_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1274" *)
  wire [12:0] _0044_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3649" *)
  wire _0045_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4509" *)
  wire _0046_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4983" *)
  wire _0047_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1412" *)
  wire [2:0] _0048_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3466" *)
  wire _0049_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4326" *)
  wire _0050_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4800" *)
  wire _0051_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3527" *)
  wire _0052_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4387" *)
  wire _0053_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4861" *)
  wire _0054_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2466" *)
  wire [7:0] _0055_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3710" *)
  wire [31:0] _0056_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4570" *)
  wire [31:0] _0057_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5044" *)
  wire [31:0] _0058_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1978" *)
  wire [6:0] _0059_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2039" *)
  wire [6:0] _0060_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3730" *)
  wire [31:0] _0061_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4590" *)
  wire [31:0] _0062_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5064" *)
  wire [31:0] _0063_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2527" *)
  wire [7:0] _0064_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3720" *)
  wire [31:0] _0065_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4580" *)
  wire [31:0] _0066_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5054" *)
  wire [31:0] _0067_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2100" *)
  wire [6:0] _0068_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2161" *)
  wire [6:0] _0069_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3740" *)
  wire [31:0] _0070_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4600" *)
  wire [31:0] _0071_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5074" *)
  wire [31:0] _0072_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1665" *)
  wire _0073_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1582" *)
  wire _0074_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3283" *)
  wire _0075_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4143" *)
  wire _0076_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4617" *)
  wire _0077_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3344" *)
  wire [2:0] _0078_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4204" *)
  wire [2:0] _0079_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4678" *)
  wire [2:0] _0080_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3405" *)
  wire _0081_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4265" *)
  wire _0082_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4739" *)
  wire _0083_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:881" *)
  wire [4:0] _0084_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:942" *)
  wire [4:0] _0085_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1003" *)
  wire [4:0] _0086_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1064" *)
  wire [4:0] _0087_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:543" *)
  wire [13:0] _0088_;
  wire [1:0] _0089_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7313" *)
  wire [12:0] _0090_;
  wire [11:0] _0091_;
  wire [13:0] _0092_;
  wire [12:0] _0093_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1807" *)
  wire _0094_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1838" *)
  wire _0095_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1838" *)
  wire _0096_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1839" *)
  wire _0097_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1839" *)
  wire _0098_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1865" *)
  wire _0099_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1865" *)
  wire _0100_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1866" *)
  wire _0101_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1953" *)
  wire _0102_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1954" *)
  wire _0103_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *)
  wire _0104_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *)
  wire _0105_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2725" *)
  wire _0106_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2728" *)
  wire _0107_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *)
  wire _0108_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *)
  wire _0109_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2759" *)
  wire _0110_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2762" *)
  wire _0111_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *)
  wire _0112_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *)
  wire _0113_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *)
  wire _0114_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3654" *)
  wire _0115_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5097" *)
  wire _0116_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5480" *)
  wire _0117_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *)
  wire _0118_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *)
  wire _0119_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *)
  wire _0120_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *)
  wire _0121_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6258" *)
  wire [511:0] _0122_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6259" *)
  wire [511:0] _0123_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6260" *)
  wire [511:0] _0124_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6261" *)
  wire [511:0] _0125_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6262" *)
  wire [511:0] _0126_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6285" *)
  wire [63:0] _0127_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6286" *)
  wire [63:0] _0128_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6287" *)
  wire [63:0] _0129_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6288" *)
  wire [63:0] _0130_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6289" *)
  wire [63:0] _0131_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6292" *)
  wire _0132_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7050" *)
  wire [511:0] _0133_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7051" *)
  wire [511:0] _0134_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7052" *)
  wire [511:0] _0135_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7053" *)
  wire [511:0] _0136_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7062" *)
  wire [511:0] _0137_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7063" *)
  wire [511:0] _0138_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7064" *)
  wire [511:0] _0139_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7065" *)
  wire [511:0] _0140_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7066" *)
  wire [511:0] _0141_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7067" *)
  wire [511:0] _0142_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7068" *)
  wire [511:0] _0143_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7069" *)
  wire [511:0] _0144_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7342" *)
  wire _0145_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7515" *)
  wire _0146_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7692" *)
  wire _0147_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7693" *)
  wire _0148_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8423" *)
  wire _0149_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7694" *)
  wire [14:0] _0150_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *)
  wire _0151_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6235" *)
  wire _0152_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6243" *)
  wire _0153_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6244" *)
  wire _0154_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6245" *)
  wire _0155_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6686" *)
  wire _0156_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1574" *)
  wire _0157_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1580" *)
  wire _0158_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1650" *)
  wire _0159_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *)
  wire _0160_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *)
  wire _0161_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *)
  wire _0162_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *)
  wire [31:0] _0163_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *)
  wire _0164_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2715" *)
  wire [31:0] _0165_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2725" *)
  wire _0166_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2728" *)
  wire _0167_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2733" *)
  wire [31:0] _0168_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *)
  wire _0169_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *)
  wire [31:0] _0170_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *)
  wire _0171_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2749" *)
  wire [31:0] _0172_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2759" *)
  wire _0173_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2762" *)
  wire _0174_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2767" *)
  wire [31:0] _0175_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:484" *)
  wire _0176_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5097" *)
  wire _0177_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5499" *)
  wire _0178_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *)
  wire _0179_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *)
  wire _0180_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *)
  wire _0181_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *)
  wire _0182_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7693" *)
  wire _0183_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1409" *)
  wire _0184_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1573" *)
  wire _0185_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1649" *)
  wire _0186_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *)
  wire _0187_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2655" *)
  wire _0188_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2667" *)
  wire _0189_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2715" *)
  wire [31:0] _0190_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2733" *)
  wire [31:0] _0191_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2749" *)
  wire [31:0] _0192_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2767" *)
  wire [31:0] _0193_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5499" *)
  wire _0194_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *)
  wire _0195_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6061" *)
  wire _0196_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6061" *)
  wire _0197_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6063" *)
  wire _0198_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6063" *)
  wire _0199_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6065" *)
  wire _0200_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6065" *)
  wire _0201_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6067" *)
  wire _0202_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6067" *)
  wire _0203_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6069" *)
  wire _0204_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6069" *)
  wire _0205_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6071" *)
  wire _0206_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6071" *)
  wire _0207_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6073" *)
  wire _0208_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6073" *)
  wire _0209_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6075" *)
  wire _0210_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6075" *)
  wire _0211_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6077" *)
  wire _0212_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6077" *)
  wire _0213_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6079" *)
  wire _0214_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6079" *)
  wire _0215_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6081" *)
  wire _0216_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6081" *)
  wire _0217_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6083" *)
  wire _0218_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6083" *)
  wire _0219_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6085" *)
  wire _0220_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6085" *)
  wire _0221_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6087" *)
  wire _0222_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6087" *)
  wire _0223_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6089" *)
  wire _0224_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6089" *)
  wire _0225_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6091" *)
  wire _0226_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6091" *)
  wire _0227_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6100" *)
  wire _0228_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6100" *)
  wire _0229_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6102" *)
  wire _0230_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6102" *)
  wire _0231_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6104" *)
  wire _0232_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6104" *)
  wire _0233_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6106" *)
  wire _0234_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6106" *)
  wire _0235_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6108" *)
  wire _0236_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6108" *)
  wire _0237_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6110" *)
  wire _0238_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6110" *)
  wire _0239_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6112" *)
  wire _0240_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6112" *)
  wire _0241_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6114" *)
  wire _0242_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6114" *)
  wire _0243_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6116" *)
  wire _0244_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6116" *)
  wire _0245_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6118" *)
  wire _0246_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6118" *)
  wire _0247_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6120" *)
  wire _0248_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6120" *)
  wire _0249_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6122" *)
  wire _0250_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6122" *)
  wire _0251_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6124" *)
  wire _0252_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6124" *)
  wire _0253_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6126" *)
  wire _0254_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6126" *)
  wire _0255_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6128" *)
  wire _0256_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6128" *)
  wire _0257_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6130" *)
  wire _0258_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6130" *)
  wire _0259_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6132" *)
  wire _0260_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6132" *)
  wire _0261_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6134" *)
  wire _0262_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6134" *)
  wire _0263_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6136" *)
  wire _0264_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6136" *)
  wire _0265_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6138" *)
  wire _0266_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6138" *)
  wire _0267_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6140" *)
  wire _0268_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6140" *)
  wire _0269_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6142" *)
  wire _0270_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6142" *)
  wire _0271_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6144" *)
  wire _0272_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6144" *)
  wire _0273_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6146" *)
  wire _0274_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6146" *)
  wire _0275_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6148" *)
  wire _0276_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6148" *)
  wire _0277_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6150" *)
  wire _0278_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6150" *)
  wire _0279_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6152" *)
  wire _0280_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6152" *)
  wire _0281_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6154" *)
  wire _0282_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6154" *)
  wire _0283_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6156" *)
  wire _0284_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6156" *)
  wire _0285_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6158" *)
  wire _0286_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6158" *)
  wire _0287_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6160" *)
  wire _0288_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6160" *)
  wire _0289_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6162" *)
  wire _0290_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6162" *)
  wire _0291_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6164" *)
  wire _0292_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6164" *)
  wire _0293_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6166" *)
  wire _0294_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6166" *)
  wire _0295_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6168" *)
  wire _0296_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6168" *)
  wire _0297_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6170" *)
  wire _0298_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6170" *)
  wire _0299_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6172" *)
  wire _0300_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6172" *)
  wire _0301_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6174" *)
  wire _0302_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6174" *)
  wire _0303_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6176" *)
  wire _0304_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6176" *)
  wire _0305_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6178" *)
  wire _0306_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6178" *)
  wire _0307_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6180" *)
  wire _0308_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6180" *)
  wire _0309_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6182" *)
  wire _0310_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6182" *)
  wire _0311_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6184" *)
  wire _0312_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6184" *)
  wire _0313_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6186" *)
  wire _0314_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6186" *)
  wire _0315_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6188" *)
  wire _0316_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6188" *)
  wire _0317_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6190" *)
  wire _0318_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6190" *)
  wire _0319_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6192" *)
  wire _0320_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6192" *)
  wire _0321_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6194" *)
  wire _0322_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6194" *)
  wire _0323_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6196" *)
  wire _0324_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6196" *)
  wire _0325_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6198" *)
  wire _0326_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6198" *)
  wire _0327_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6200" *)
  wire _0328_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6200" *)
  wire _0329_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6202" *)
  wire _0330_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6202" *)
  wire _0331_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6204" *)
  wire _0332_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6204" *)
  wire _0333_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6206" *)
  wire _0334_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6206" *)
  wire _0335_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6208" *)
  wire _0336_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6208" *)
  wire _0337_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6210" *)
  wire _0338_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6210" *)
  wire _0339_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6212" *)
  wire _0340_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6212" *)
  wire _0341_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6214" *)
  wire _0342_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6214" *)
  wire _0343_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6216" *)
  wire _0344_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6216" *)
  wire _0345_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6218" *)
  wire _0346_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6218" *)
  wire _0347_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6220" *)
  wire _0348_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6220" *)
  wire _0349_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6222" *)
  wire _0350_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6222" *)
  wire _0351_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6224" *)
  wire _0352_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6224" *)
  wire _0353_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6226" *)
  wire _0354_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6226" *)
  wire _0355_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6259" *)
  wire [511:0] _0356_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6260" *)
  wire [511:0] _0357_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6261" *)
  wire [511:0] _0358_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6286" *)
  wire [63:0] _0359_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6287" *)
  wire [63:0] _0360_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6288" *)
  wire [63:0] _0361_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *)
  wire _0362_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7051" *)
  wire [511:0] _0363_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7052" *)
  wire [511:0] _0364_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7063" *)
  wire [511:0] _0365_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7064" *)
  wire [511:0] _0366_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7065" *)
  wire [511:0] _0367_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7066" *)
  wire [511:0] _0368_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7067" *)
  wire [511:0] _0369_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7068" *)
  wire [511:0] _0370_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7507" *)
  wire _0371_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7692" *)
  wire _0372_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1259" *)
  wire _0373_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6817" *)
  wire _0374_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *)
  wire _0375_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *)
  wire [31:0] _0376_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *)
  wire [31:0] _0377_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2714" *)
  wire [31:0] _0378_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *)
  wire [31:0] _0379_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *)
  wire [31:0] _0380_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2748" *)
  wire [31:0] _0381_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1743" *)
  wire _0382_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1743" *)
  wire _0383_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2684" *)
  wire [13:0] _0384_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2699" *)
  wire [13:0] _0385_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2710" *)
  wire [31:0] _0386_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2713" *)
  wire [31:0] _0387_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2726" *)
  wire [31:0] _0388_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2729" *)
  wire [31:0] _0389_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2732" *)
  wire [31:0] _0390_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2744" *)
  wire [31:0] _0391_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2747" *)
  wire [31:0] _0392_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2760" *)
  wire [31:0] _0393_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2763" *)
  wire [31:0] _0394_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2766" *)
  wire [31:0] _0395_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7293" *)
  wire [11:0] _0396_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7304" *)
  wire [3:0] _0397_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7680" *)
  wire [2:0] _0398_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8424" *)
  wire _0399_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:116" *)
  wire [1535:0] dat_16b_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:117" *)
  wire [1535:0] dat_8b_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:118" *)
  wire [511:0] dat_l0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:119" *)
  wire [1023:0] dat_l1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:120" *)
  wire [511:0] dat_l1_hi;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:121" *)
  wire [511:0] dat_l1_lo;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:122" *)
  wire [1535:0] dat_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:204" *)
  reg [5:0] data_planar0_add;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:205" *)
  wire [5:0] data_planar0_add_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:206" *)
  reg [13:0] data_planar0_cur_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:207" *)
  wire [13:0] data_planar0_cur_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:208" *)
  wire data_planar0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:210" *)
  wire data_planar0_ori_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:211" *)
  wire [13:0] data_planar0_p0_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:212" *)
  wire [2:0] data_planar0_p0_cur_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:213" *)
  wire [31:0] data_planar0_p0_lp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:214" *)
  wire [31:0] data_planar0_p0_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:215" *)
  wire [31:0] data_planar0_p0_rp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:216" *)
  wire [31:0] data_planar0_p0_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:217" *)
  wire [13:0] data_planar0_p1_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:218" *)
  wire [2:0] data_planar0_p1_cur_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:219" *)
  reg [2:0] data_planar0_p1_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:220" *)
  wire [2:0] data_planar0_p1_flag_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:221" *)
  wire [31:0] data_planar0_p1_lp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:223" *)
  wire [31:0] data_planar0_p1_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:224" *)
  wire [31:0] data_planar0_p1_rp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:225" *)
  wire [31:0] data_planar0_p1_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:226" *)
  reg [5:0] data_planar1_add;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:227" *)
  wire [5:0] data_planar1_add_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:228" *)
  reg [13:0] data_planar1_cur_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:229" *)
  wire [13:0] data_planar1_cur_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:230" *)
  wire data_planar1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:232" *)
  wire data_planar1_ori_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:233" *)
  wire [13:0] data_planar1_p0_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:234" *)
  wire [2:0] data_planar1_p0_cur_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:235" *)
  wire [31:0] data_planar1_p0_lp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:236" *)
  wire [31:0] data_planar1_p0_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:237" *)
  wire [31:0] data_planar1_p0_rp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:238" *)
  wire [31:0] data_planar1_p0_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:239" *)
  wire [13:0] data_planar1_p1_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:240" *)
  wire [2:0] data_planar1_p1_cur_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:241" *)
  reg [2:0] data_planar1_p1_flag;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:242" *)
  wire [2:0] data_planar1_p1_flag_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:243" *)
  wire [31:0] data_planar1_p1_lp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:245" *)
  wire [31:0] data_planar1_p1_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:246" *)
  wire [31:0] data_planar1_p1_rp_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:247" *)
  wire [31:0] data_planar1_p1_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:123" *)
  wire [13:0] data_width_mark_0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:248" *)
  reg [13:0] data_width_mark_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:124" *)
  wire [13:0] data_width_mark_1_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:249" *)
  reg [13:0] data_width_mark_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:125" *)
  wire [13:0] data_width_mark_2_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:91" *)
  output [11:0] img2cvt_dat_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:92" *)
  output [1023:0] img2cvt_dat_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:93" *)
  output img2cvt_dat_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:94" *)
  output img2cvt_dat_wr_hsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:95" *)
  output [11:0] img2cvt_dat_wr_info_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:115" *)
  output [127:0] img2cvt_dat_wr_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:96" *)
  output [1023:0] img2cvt_mn_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:97" *)
  output [7:0] img2sbuf_p0_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:65" *)
  input [255:0] img2sbuf_p0_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:98" *)
  output img2sbuf_p0_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:99" *)
  output [7:0] img2sbuf_p1_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:66" *)
  input [255:0] img2sbuf_p1_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:100" *)
  output img2sbuf_p1_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:101" *)
  output [11:0] img2status_dat_entries;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:102" *)
  output [11:0] img2status_dat_slices;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:103" *)
  output img2status_dat_updt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:126" *)
  wire img_layer_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:127" *)
  wire img_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:128" *)
  wire [3:0] img_p0_burst;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:129" *)
  (* unused_bits = "1 2 3 4" *)
  wire [4:0] img_p1_burst;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:130" *)
  (* unused_bits = "5 6 7 8" *)
  wire [10:0] img_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:250" *)
  wire is_1st_height;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:251" *)
  wire is_addr_wrap;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:252" *)
  wire is_base_wrap;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:253" *)
  wire is_first_running;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:254" *)
  wire is_last_height;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:255" *)
  wire is_last_loop;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:256" *)
  wire is_last_pburst;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:257" *)
  wire is_last_planar;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:131" *)
  wire is_last_sub_h;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:67" *)
  input is_running;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:258" *)
  reg is_running_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:68" *)
  input layer_st;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:259" *)
  reg [4:0] lp_planar0_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:260" *)
  wire [4:0] lp_planar0_mask_sft_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:261" *)
  reg [4:0] lp_planar1_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:262" *)
  wire [4:0] lp_planar1_mask_sft_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:132" *)
  wire [63:0] mask_pad;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:263" *)
  reg [63:0] mask_pad_planar0_c0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:264" *)
  reg [63:0] mask_pad_planar1_c0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:265" *)
  reg [63:0] mask_pad_planar1_c1_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:133" *)
  wire [63:0] mask_zero;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:266" *)
  wire [511:0] mn_16b_mnorm;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:267" *)
  wire [1535:0] mn_16b_myuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:268" *)
  wire [1023:0] mn_8b_mnorm;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:269" *)
  wire [3071:0] mn_8b_myuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:134" *)
  wire [1023:0] mn_ch1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:135" *)
  wire [1023:0] mn_ch1_4;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:136" *)
  wire [3071:0] mn_ch3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:137" *)
  wire [1023:0] mn_ch4;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:138" *)
  (* unused_bits = "64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127" *)
  wire [127:0] mn_mask_uv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:139" *)
  wire mn_mask_uv_0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:140" *)
  wire mn_mask_uv_1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:141" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" *)
  wire [63:0] mn_mask_uv_hi;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:142" *)
  wire [63:0] mn_mask_uv_lo;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:271" *)
  reg [63:0] mn_mask_uv_lo_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:143" *)
  wire [63:0] mn_mask_y;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:272" *)
  reg [63:0] mn_mask_y_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:144" *)
  wire mn_mask_y_en;
  (* unused_bits = "98 99 100 101 104 105 106 107 110 111 112 113 116 117 118 119 122 123 124 125 128 129 130 131 134 135 136 137 140 141 142 143 146 147 148 149 152 153 154 155 158 159 160 161 164 165 166 167 170 171 172 173 176 177 178 179 182 183 184 185" *)
  wire [187:0] mn_mask_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:281" *)
  wire mon_pk_rsp_wr_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:282" *)
  wire mon_pk_rsp_wr_h_offset_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:283" *)
  wire mon_pk_rsp_wr_w_offset_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:63" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:64" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:104" *)
  output pack_is_done;
  reg pack_is_done;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:291" *)
  wire pack_is_done_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:292" *)
  reg [4:0] pad_left_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:146" *)
  wire [191:0] pad_mask_16b_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:147" *)
  wire [191:0] pad_mask_8b_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:148" *)
  wire [63:0] pad_mask_l0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:149" *)
  wire [127:0] pad_mask_l1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:150" *)
  wire [63:0] pad_mask_l1_hi;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:151" *)
  wire [63:0] pad_mask_l1_lo;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:152" *)
  wire [191:0] pad_mask_yuv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:69" *)
  input [3:0] pixel_bank;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:70" *)
  input pixel_data_expand;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:71" *)
  input pixel_data_shrink;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:72" *)
  input pixel_early_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:73" *)
  input pixel_packed_10b;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:74" *)
  input pixel_planar;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:75" *)
  input [2:0] pixel_planar0_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:76" *)
  input [2:0] pixel_planar1_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:77" *)
  input [1:0] pixel_precision;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:78" *)
  input pixel_uint;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:153" *)
  wire [1023:0] pk_mn_out_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:293" *)
  reg [511:0] pk_mn_out_data_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:294" *)
  reg [511:0] pk_mn_out_data_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:295" *)
  reg [11:0] pk_out_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:154" *)
  wire [1023:0] pk_out_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:296" *)
  reg [11:0] pk_out_data_entries;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:297" *)
  reg [511:0] pk_out_data_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:298" *)
  reg [511:0] pk_out_data_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:299" *)
  reg [3:0] pk_out_data_slices;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:300" *)
  reg pk_out_data_updt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:301" *)
  reg pk_out_ext128;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:302" *)
  reg pk_out_ext64;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:303" *)
  reg pk_out_hsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:155" *)
  wire [11:0] pk_out_info_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:156" *)
  wire pk_out_interleave;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:304" *)
  reg [3:0] pk_out_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:305" *)
  reg pk_out_mean;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:157" *)
  wire [127:0] pk_out_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:306" *)
  reg [63:0] pk_out_pad_mask_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:307" *)
  reg [63:0] pk_out_pad_mask_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:308" *)
  reg [2:0] pk_out_sub_h;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:309" *)
  reg pk_out_uint;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:310" *)
  reg pk_out_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:158" *)
  wire pk_rsp_1st_height;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:311" *)
  reg pk_rsp_1st_height_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:159" *)
  wire pk_rsp_cur_1st_height;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:160" *)
  wire pk_rsp_cur_layer_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:161" *)
  wire pk_rsp_cur_loop_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:162" *)
  wire pk_rsp_cur_one_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:163" *)
  wire [2:0] pk_rsp_cur_sub_h;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:164" *)
  wire pk_rsp_cur_sub_h_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:165" *)
  wire pk_rsp_cur_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:166" *)
  wire [1023:0] pk_rsp_dat_ergb;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:312" *)
  wire [1023:0] pk_rsp_dat_mergb;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:313" *)
  wire [511:0] pk_rsp_dat_mnorm;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:167" *)
  wire [511:0] pk_rsp_dat_normal;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:168" *)
  wire [11:0] pk_rsp_data_entries;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:314" *)
  wire [511:0] pk_rsp_data_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:169" *)
  wire pk_rsp_data_h0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:315" *)
  wire [511:0] pk_rsp_data_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:170" *)
  wire pk_rsp_data_h1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:171" *)
  wire [3:0] pk_rsp_data_slices;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:316" *)
  wire pk_rsp_data_updt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:172" *)
  wire pk_rsp_early_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:173" *)
  wire pk_rsp_layer_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:317" *)
  reg pk_rsp_layer_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:174" *)
  wire pk_rsp_loop_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:318" *)
  reg pk_rsp_loop_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:319" *)
  wire [511:0] pk_rsp_mn_data_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:175" *)
  wire pk_rsp_mn_data_h0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:320" *)
  wire [511:0] pk_rsp_mn_data_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:176" *)
  wire pk_rsp_mn_data_h1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:321" *)
  wire [7:0] pk_rsp_mn_sel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:177" *)
  wire pk_rsp_one_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:322" *)
  reg pk_rsp_one_line_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:323" *)
  wire [4:0] pk_rsp_out_sel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:178" *)
  wire [255:0] pk_rsp_p0_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:179" *)
  wire [31:0] pk_rsp_p0_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:180" *)
  wire [31:0] pk_rsp_p0_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:181" *)
  wire [255:0] pk_rsp_p1_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:182" *)
  wire [31:0] pk_rsp_p1_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:183" *)
  wire [31:0] pk_rsp_p1_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:184" *)
  wire [127:0] pk_rsp_pad_mask_ergb;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:324" *)
  wire [63:0] pk_rsp_pad_mask_h0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:325" *)
  wire [63:0] pk_rsp_pad_mask_h1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:185" *)
  wire [63:0] pk_rsp_pad_mask_norm;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:186" *)
  wire pk_rsp_pipe_sel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:187" *)
  wire pk_rsp_planar;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:326" *)
  reg [511:0] pk_rsp_planar0_c0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:188" *)
  wire pk_rsp_planar0_c0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:327" *)
  reg [511:0] pk_rsp_planar1_c0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:189" *)
  wire pk_rsp_planar1_c0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:328" *)
  reg [511:0] pk_rsp_planar1_c1_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:190" *)
  wire pk_rsp_planar1_c1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:191" *)
  wire [2:0] pk_rsp_sub_h;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:329" *)
  reg [2:0] pk_rsp_sub_h_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:192" *)
  wire pk_rsp_sub_h_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:330" *)
  reg pk_rsp_sub_h_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:193" *)
  wire pk_rsp_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:331" *)
  reg pk_rsp_vld_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:194" *)
  wire pk_rsp_vld_d1_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:332" *)
  wire [11:0] pk_rsp_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:333" *)
  wire [13:0] pk_rsp_wr_addr_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:334" *)
  wire [3:0] pk_rsp_wr_addr_wrap;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:335" *)
  reg [11:0] pk_rsp_wr_base;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:336" *)
  wire pk_rsp_wr_base_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:337" *)
  wire [12:0] pk_rsp_wr_base_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:338" *)
  wire [11:0] pk_rsp_wr_base_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:339" *)
  wire [3:0] pk_rsp_wr_base_wrap;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:340" *)
  reg [1:0] pk_rsp_wr_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:341" *)
  wire [1:0] pk_rsp_wr_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:342" *)
  wire [11:0] pk_rsp_wr_entries;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:195" *)
  wire pk_rsp_wr_ext128;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:196" *)
  wire pk_rsp_wr_ext64;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:343" *)
  reg [11:0] pk_rsp_wr_h_offset;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:344" *)
  wire pk_rsp_wr_h_offset_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:345" *)
  wire [11:0] pk_rsp_wr_h_offset_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:197" *)
  wire [3:0] pk_rsp_wr_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:198" *)
  wire [2:0] pk_rsp_wr_size_ori;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:346" *)
  wire [3:0] pk_rsp_wr_slices;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:199" *)
  wire [1:0] pk_rsp_wr_sub_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:347" *)
  wire pk_rsp_wr_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:348" *)
  wire [2:0] pk_rsp_wr_w_add;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:349" *)
  reg [13:0] pk_rsp_wr_w_offset;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:350" *)
  wire pk_rsp_wr_w_offset_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:351" *)
  reg [13:0] pk_rsp_wr_w_offset_ori;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:352" *)
  wire pk_rsp_wr_w_offset_ori_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:353" *)
  wire [13:0] pk_rsp_wr_w_offset_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:354" *)
  reg rd_1st_height_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:355" *)
  reg rd_1st_height_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:356" *)
  reg rd_1st_height_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:357" *)
  reg [12:0] rd_height_cnt;
  wire [12:0] rd_height_cnt_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:359" *)
  wire [12:0] rd_height_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:360" *)
  wire rd_height_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:361" *)
  wire rd_height_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:362" *)
  wire [1:0] rd_idx_add;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:363" *)
  reg rd_layer_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:364" *)
  reg rd_layer_end_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:365" *)
  reg rd_layer_end_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:366" *)
  wire rd_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:367" *)
  reg rd_local_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:368" *)
  wire rd_local_vld_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:369" *)
  reg [2:0] rd_loop_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:370" *)
  wire [2:0] rd_loop_cnt_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:371" *)
  wire [2:0] rd_loop_cnt_limit;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:372" *)
  wire [2:0] rd_loop_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:373" *)
  wire rd_loop_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:374" *)
  wire rd_loop_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:375" *)
  reg rd_loop_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:376" *)
  reg rd_loop_end_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:377" *)
  reg rd_loop_end_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:378" *)
  reg rd_one_line_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:379" *)
  reg rd_one_line_end_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:380" *)
  reg rd_one_line_end_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:381" *)
  wire [7:0] rd_p0_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:382" *)
  reg [7:0] rd_p0_addr_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:383" *)
  wire [31:0] rd_p0_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:384" *)
  reg [31:0] rd_p0_pad_mask_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:385" *)
  reg [31:0] rd_p0_pad_mask_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:386" *)
  reg [31:0] rd_p0_pad_mask_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:387" *)
  reg [6:0] rd_p0_planar0_idx;
  wire [6:0] rd_p0_planar0_idx_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:389" *)
  wire [6:0] rd_p0_planar0_idx_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:391" *)
  reg [6:0] rd_p0_planar1_idx;
  wire [6:0] rd_p0_planar1_idx_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:393" *)
  wire [6:0] rd_p0_planar1_idx_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:395" *)
  wire rd_p0_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:396" *)
  reg rd_p0_vld_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:397" *)
  wire [31:0] rd_p0_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:398" *)
  reg [31:0] rd_p0_zero_mask_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:399" *)
  reg [31:0] rd_p0_zero_mask_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:400" *)
  reg [31:0] rd_p0_zero_mask_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:401" *)
  wire [7:0] rd_p1_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:402" *)
  reg [7:0] rd_p1_addr_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:403" *)
  wire [31:0] rd_p1_pad_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:404" *)
  reg [31:0] rd_p1_pad_mask_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:405" *)
  reg [31:0] rd_p1_pad_mask_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:406" *)
  reg [31:0] rd_p1_pad_mask_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:407" *)
  reg [6:0] rd_p1_planar0_idx;
  wire [6:0] rd_p1_planar0_idx_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:409" *)
  wire [6:0] rd_p1_planar0_idx_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:411" *)
  reg [6:0] rd_p1_planar1_idx;
  wire [6:0] rd_p1_planar1_idx_inc;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:413" *)
  wire [6:0] rd_p1_planar1_idx_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:415" *)
  wire rd_p1_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:416" *)
  reg rd_p1_vld_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:417" *)
  wire [31:0] rd_p1_zero_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:418" *)
  reg [31:0] rd_p1_zero_mask_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:419" *)
  reg [31:0] rd_p1_zero_mask_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:420" *)
  reg [31:0] rd_p1_zero_mask_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:421" *)
  reg rd_pburst_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:422" *)
  wire rd_pburst_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:423" *)
  wire rd_pburst_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:424" *)
  wire rd_pburst_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:425" *)
  wire rd_pburst_limit;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:427" *)
  wire rd_planar0_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:428" *)
  wire rd_planar0_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:429" *)
  wire rd_planar0_ori_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:430" *)
  wire [1:0] rd_planar0_rd_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:432" *)
  wire rd_planar1_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:433" *)
  wire rd_planar1_line_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:434" *)
  wire rd_planar1_ori_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:435" *)
  wire [1:0] rd_planar1_rd_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:436" *)
  reg rd_planar_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:437" *)
  wire rd_planar_cnt_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:438" *)
  reg rd_planar_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:439" *)
  reg rd_planar_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:440" *)
  reg rd_planar_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:441" *)
  wire rd_planar_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:442" *)
  wire rd_planar_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:443" *)
  wire [1:0] rd_rd_mask;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:200" *)
  wire [2:0] rd_sub_h_cnt;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:444" *)
  reg [2:0] rd_sub_h_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:445" *)
  reg [2:0] rd_sub_h_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:446" *)
  reg [2:0] rd_sub_h_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:447" *)
  wire rd_sub_h_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:448" *)
  reg rd_sub_h_end_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:449" *)
  reg rd_sub_h_end_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:450" *)
  reg rd_sub_h_end_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:451" *)
  wire rd_vld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:452" *)
  reg rd_vld_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:453" *)
  reg rd_vld_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:454" *)
  reg rd_vld_d3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:201" *)
  wire [511:0] rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:107" *)
  input [12:0] reg2dp_datain_channel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:106" *)
  input [12:0] reg2dp_datain_width;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:111" *)
  input [15:0] reg2dp_mean_ax;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:110" *)
  input [15:0] reg2dp_mean_bv;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:109" *)
  input [15:0] reg2dp_mean_gu;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:108" *)
  input [15:0] reg2dp_mean_ry;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:112" *)
  input [4:0] reg2dp_pad_left;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:113" *)
  input [5:0] reg2dp_pad_right;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:455" *)
  reg [4:0] rp_planar0_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:456" *)
  wire [4:0] rp_planar0_mask_sft_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:457" *)
  reg [4:0] rp_planar1_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:458" *)
  wire [4:0] rp_planar1_mask_sft_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:79" *)
  input [11:0] sg2pack_data_entries;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:80" *)
  input [11:0] sg2pack_entry_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:81" *)
  input [11:0] sg2pack_entry_mid;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:82" *)
  input [11:0] sg2pack_entry_st;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:83" *)
  input [12:0] sg2pack_height_total;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:84" *)
  input [10:0] sg2pack_img_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:105" *)
  output sg2pack_img_prdy;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:85" *)
  input sg2pack_img_pvld;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:86" *)
  input sg2pack_mn_enable;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:87" *)
  input [3:0] sg2pack_sub_h_end;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:88" *)
  input [3:0] sg2pack_sub_h_mid;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:89" *)
  input [3:0] sg2pack_sub_h_st;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:90" *)
  input [11:0] status2dma_wr_idx;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:202" *)
  wire [13:0] z14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:203" *)
  wire [5:0] z6;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:459" *)
  reg [4:0] zero_planar0_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:460" *)
  wire [4:0] zero_planar0_mask_sft_w;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:461" *)
  reg [4:0] zero_planar1_mask_sft;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:462" *)
  wire [4:0] zero_planar1_mask_sft_w;
  assign rd_height_cnt_inc = rd_height_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1254" *) 1'b1;
  assign rd_loop_cnt_limit = img_pd[3:1] + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1390" *) img_pd[0];
  assign rd_loop_cnt_inc = rd_loop_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1396" *) 1'b1;
  assign rd_p0_planar0_idx_inc = rd_p0_planar0_idx + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1909" *) rd_idx_add;
  assign rd_p1_planar0_idx_inc = rd_p1_planar0_idx + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1910" *) rd_idx_add;
  assign rd_p0_planar1_idx_inc = rd_p0_planar1_idx + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1911" *) rd_idx_add;
  assign rd_p1_planar1_idx_inc = rd_p1_planar1_idx + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1912" *) rd_idx_add;
  assign data_planar0_p0_cnt_w = data_planar0_cur_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2594" *) data_planar0_add;
  assign data_planar0_p1_cnt_w = data_planar0_cur_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2596" *) { data_planar0_add, 1'b0 };
  assign data_planar1_p0_cnt_w = data_planar1_cur_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2603" *) data_planar1_add;
  assign data_planar1_p1_cnt_w = data_planar1_cur_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2605" *) { data_planar1_add, 1'b0 };
  assign _0088_ = reg2dp_pad_left + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:543" *) reg2dp_datain_width;
  assign data_width_mark_1_w = _0088_ + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:543" *) 1'b1;
  assign data_width_mark_2_w = data_width_mark_1_w + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:544" *) reg2dp_pad_right;
  assign _0089_ = pk_rsp_wr_cnt + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5500" *) 1'b1;
  assign _0090_ = pk_rsp_wr_base + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7313" *) pk_rsp_data_entries;
  assign _0091_ = pk_rsp_wr_h_offset + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7508" *) sg2pack_data_entries;
  assign _0092_ = pk_rsp_wr_w_offset + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7694" *) pk_rsp_wr_w_add;
  assign _0093_ = pk_rsp_wr_base + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7972" *) pk_rsp_wr_h_offset;
  assign pk_rsp_wr_addr_inc = _0093_ + (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7972" *) pk_rsp_wr_w_offset[13:2];
  assign rd_pburst_limit = rd_planar_cnt & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *) _0187_;
  assign sg2pack_img_prdy = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1727" *) rd_loop_end;
  assign rd_pburst_end = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1749" *) is_last_pburst;
  assign rd_planar_end = rd_pburst_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1756" *) is_last_planar;
  assign rd_loop_end = rd_planar_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1764" *) is_last_loop;
  assign rd_line_end = rd_loop_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1783" *) img_pd[9];
  assign rd_height_end = rd_line_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1794" *) is_last_height;
  assign _0094_ = rd_pburst_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1807" *) pixel_planar;
  assign _0095_ = rd_pburst_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1838" *) _0157_;
  assign _0096_ = _0095_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1838" *) is_last_loop;
  assign rd_planar0_line_end = _0096_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1838" *) img_pd[9];
  assign _0097_ = rd_pburst_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1839" *) rd_planar_cnt;
  assign _0098_ = _0097_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1839" *) is_last_loop;
  assign rd_planar1_line_end = _0098_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1839" *) img_pd[9];
  assign _0099_ = is_last_loop & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1865" *) is_last_pburst;
  assign _0100_ = _0099_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1865" *) img_pd[0];
  assign _0101_ = _0099_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1866" *) img_pd[4];
  assign rd_p0_vld = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1879" *) rd_rd_mask[0];
  assign rd_p1_vld = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1880" *) rd_rd_mask[1];
  assign _0102_ = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1953" *) _0157_;
  assign _0103_ = rd_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1954" *) rd_planar_cnt;
  assign _0104_ = _0162_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *) data_planar0_p0_cur_flag[0];
  assign _0105_ = _0164_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *) data_planar0_p0_cur_flag[1];
  assign data_planar0_p0_pad_mask = _0190_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2715" *) _0165_;
  assign _0106_ = _0166_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2725" *) data_planar0_p1_cur_flag[0];
  assign _0107_ = _0167_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2728" *) data_planar0_p1_cur_flag[1];
  assign data_planar0_p1_pad_mask = _0191_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2733" *) _0168_;
  assign _0108_ = _0169_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *) data_planar1_p0_cur_flag[0];
  assign _0109_ = _0171_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *) data_planar1_p0_cur_flag[1];
  assign data_planar1_p0_pad_mask = _0192_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2749" *) _0172_;
  assign _0110_ = _0173_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2759" *) data_planar1_p1_cur_flag[0];
  assign _0111_ = _0174_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2762" *) data_planar1_p1_cur_flag[1];
  assign data_planar1_p1_pad_mask = _0193_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2767" *) _0175_;
  assign _0112_ = is_last_pburst & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *) is_last_planar;
  assign _0113_ = _0112_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *) is_last_loop;
  assign _0114_ = _0113_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3532" *) img_pd[9];
  assign _0115_ = img_pd[10] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3654" *) rd_height_end;
  assign is_first_running = _0176_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:484" *) is_running;
  assign pk_rsp_early_end = pixel_early_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5096" *) rd_one_line_end_d3;
  assign _0116_ = rd_vld_d3 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5097" *) pixel_planar;
  assign pk_rsp_vld_d1_w = _0116_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5097" *) _0177_;
  assign _0117_ = rd_vld_d3 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5480" *) pk_rsp_early_end;
  assign _0118_ = pk_rsp_cur_one_line_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *) _0151_;
  assign _0119_ = _0118_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *) pixel_data_shrink;
  assign pk_rsp_wr_ext64 = _0119_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *) _0179_;
  assign _0120_ = pk_rsp_cur_one_line_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) _0180_;
  assign _0121_ = _0181_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) _0179_;
  assign pk_rsp_wr_ext128 = _0120_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) _0195_;
  assign pk_rsp_out_sel[1] = _0158_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6242" *) _0179_;
  assign pk_rsp_out_sel[2] = pixel_planar & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6243" *) _0153_;
  assign pk_rsp_out_sel[3] = pixel_planar & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6244" *) _0154_;
  assign pk_rsp_out_sel[4] = pixel_planar & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6245" *) _0155_;
  assign _0122_ = { pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6258" *) pk_rsp_dat_mergb[511:0];
  assign _0123_ = { pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6259" *) pk_rsp_dat_mnorm;
  assign _0124_ = { pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6260" *) dat_yuv[511:0];
  assign _0125_ = { pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6261" *) dat_yuv[1023:512];
  assign _0126_ = { pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6262" *) { dat_l1_hi[511:496], dat_yuv[1519:1024] };
  assign _0127_ = { pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b, pixel_packed_10b } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6285" *) { rd_p0_pad_mask_d3[31], rd_p0_pad_mask_d3[31:30], rd_p0_pad_mask_d3[30:29], rd_p0_pad_mask_d3[29:28], rd_p0_pad_mask_d3[28:27], rd_p0_pad_mask_d3[27:26], rd_p0_pad_mask_d3[26:25], rd_p0_pad_mask_d3[25:24], rd_p0_pad_mask_d3[24:23], rd_p0_pad_mask_d3[23:22], rd_p0_pad_mask_d3[22:21], rd_p0_pad_mask_d3[21:20], rd_p0_pad_mask_d3[20:19], rd_p0_pad_mask_d3[19:18], rd_p0_pad_mask_d3[18:17], rd_p0_pad_mask_d3[17:16], rd_p0_pad_mask_d3[16:15], rd_p0_pad_mask_d3[15:14], rd_p0_pad_mask_d3[14:13], rd_p0_pad_mask_d3[13:12], rd_p0_pad_mask_d3[12:11], rd_p0_pad_mask_d3[11:10], rd_p0_pad_mask_d3[10:9], rd_p0_pad_mask_d3[9:8], rd_p0_pad_mask_d3[8:7], rd_p0_pad_mask_d3[7:6], rd_p0_pad_mask_d3[6:5], rd_p0_pad_mask_d3[5:4], rd_p0_pad_mask_d3[4:3], rd_p0_pad_mask_d3[3:2], rd_p0_pad_mask_d3[2:1], rd_p0_pad_mask_d3[1:0], rd_p0_pad_mask_d3[0] };
  assign _0128_ = { pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1], pk_rsp_out_sel[1] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6286" *) { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 };
  assign _0129_ = { pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2], pk_rsp_out_sel[2] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6287" *) pad_mask_yuv[63:0];
  assign _0130_ = { pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3], pk_rsp_out_sel[3] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6288" *) pad_mask_yuv[127:64];
  assign _0131_ = { pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4], pk_rsp_out_sel[4] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6289" *) { pad_mask_l1_hi[63:62], pad_mask_yuv[189:128] };
  assign mn_mask_y_en = _0116_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6291" *) _0178_;
  assign _0132_ = _0116_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6292" *) rd_planar_d3;
  assign mn_mask_uv_0_en = _0132_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6292" *) _0153_;
  assign pk_rsp_planar1_c1_en = _0132_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6293" *) _0154_;
  assign pk_rsp_data_h1_en = pk_rsp_wr_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6295" *) pixel_packed_10b;
  assign pk_rsp_mn_sel[0] = _0158_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *) _0362_;
  assign pk_rsp_mn_sel[1] = pk_rsp_out_sel[1] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7037" *) _0375_;
  assign pk_rsp_mn_sel[2] = pk_rsp_out_sel[2] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7038" *) _0182_;
  assign pk_rsp_mn_sel[3] = pk_rsp_out_sel[2] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7039" *) _0375_;
  assign pk_rsp_mn_sel[4] = pk_rsp_out_sel[3] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7040" *) _0182_;
  assign pk_rsp_mn_sel[5] = pk_rsp_out_sel[3] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7041" *) _0375_;
  assign pk_rsp_mn_sel[6] = pk_rsp_out_sel[4] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7042" *) _0182_;
  assign pk_rsp_mn_sel[7] = pk_rsp_out_sel[4] & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7043" *) _0375_;
  assign _0133_ = { pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7050" *) mn_8b_mnorm[1023:512];
  assign _0134_ = { pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7051" *) { mn_8b_myuv[1023:1008], mn_16b_myuv[527:480], mn_8b_myuv[959:912], mn_16b_myuv[479:432], mn_8b_myuv[863:816], mn_16b_myuv[431:384], mn_8b_myuv[767:720], mn_16b_myuv[383:336], mn_8b_myuv[671:624], mn_16b_myuv[335:288], mn_8b_myuv[575:528], mn_16b_myuv[287:272] };
  assign _0135_ = { pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7052" *) { mn_16b_myuv[1039:1008], mn_8b_myuv[2015:1968], mn_16b_myuv[1007:960], mn_8b_myuv[1919:1872], mn_16b_myuv[959:912], mn_8b_myuv[1823:1776], mn_16b_myuv[911:864], mn_8b_myuv[1727:1680], mn_16b_myuv[863:816], mn_8b_myuv[1631:1584], mn_16b_myuv[815:768] };
  assign _0136_ = { pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7053" *) { mn_8b_myuv[3071:3024], mn_16b_myuv[1535:1488], mn_8b_myuv[2975:2928], mn_16b_myuv[1487:1440], mn_8b_myuv[2879:2832], mn_16b_myuv[1439:1392], mn_8b_myuv[2783:2736], mn_16b_myuv[1391:1344], mn_8b_myuv[2687:2640], mn_16b_myuv[1343:1296], mn_8b_myuv[2591:2560] };
  assign _0137_ = { pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0], pk_rsp_mn_sel[0] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7062" *) { mn_8b_mnorm[511:16], mn_16b_mnorm[15:0] };
  assign _0138_ = { pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1], pk_rsp_mn_sel[1] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7063" *) mn_16b_mnorm;
  assign _0139_ = { pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2], pk_rsp_mn_sel[2] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7064" *) { mn_16b_myuv[271:240], mn_8b_myuv[479:432], mn_16b_myuv[239:192], mn_8b_myuv[383:336], mn_16b_myuv[191:144], mn_8b_myuv[287:240], mn_16b_myuv[143:96], mn_8b_myuv[191:144], mn_16b_myuv[95:48], mn_8b_myuv[95:48], mn_16b_myuv[47:0] };
  assign _0140_ = { pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3], pk_rsp_mn_sel[3] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7065" *) mn_16b_myuv[511:0];
  assign _0141_ = { pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4], pk_rsp_mn_sel[4] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7066" *) { mn_8b_myuv[1535:1488], mn_16b_myuv[767:720], mn_8b_myuv[1439:1392], mn_16b_myuv[719:672], mn_8b_myuv[1343:1296], mn_16b_myuv[671:624], mn_8b_myuv[1247:1200], mn_16b_myuv[623:576], mn_8b_myuv[1151:1104], mn_16b_myuv[575:528], mn_8b_myuv[1055:1024] };
  assign _0142_ = { pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5], pk_rsp_mn_sel[5] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7067" *) mn_16b_myuv[1023:512];
  assign _0143_ = { pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6], pk_rsp_mn_sel[6] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7068" *) { mn_8b_myuv[2559:2544], mn_16b_myuv[1295:1248], mn_8b_myuv[2495:2448], mn_16b_myuv[1247:1200], mn_8b_myuv[2399:2352], mn_16b_myuv[1199:1152], mn_8b_myuv[2303:2256], mn_16b_myuv[1151:1104], mn_8b_myuv[2207:2160], mn_16b_myuv[1103:1056], mn_8b_myuv[2111:2064], mn_16b_myuv[1055:1040] };
  assign _0144_ = { pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7], pk_rsp_mn_sel[7] } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7069" *) mn_16b_myuv[1535:1024];
  assign pk_rsp_mn_data_h1_en = pk_rsp_wr_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7075" *) _0362_;
  assign _0145_ = pk_rsp_wr_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7342" *) pk_rsp_cur_one_line_end;
  assign pk_rsp_data_updt = _0145_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7342" *) pk_rsp_cur_sub_h_end;
  assign _0146_ = pk_rsp_wr_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7515" *) pk_rsp_cur_loop_end;
  assign _0147_ = pk_rsp_cur_one_line_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7692" *) pk_rsp_cur_sub_h_end;
  assign _0148_ = pk_rsp_cur_loop_end & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7693" *) _0183_;
  assign _0149_ = pk_rsp_wr_vld & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8423" *) pk_rsp_cur_layer_end;
  assign is_last_height = rd_height_cnt == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1265" *) sg2pack_height_total;
  assign is_last_pburst = rd_pburst_cnt == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1663" *) rd_pburst_limit;
  assign _0151_ = pk_rsp_wr_w_offset[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *) 2'b10;
  assign _0152_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6235" *) pixel_precision;
  assign _0153_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6243" *) pk_rsp_wr_cnt;
  assign _0154_ = pk_rsp_wr_cnt == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6244" *) 1'b1;
  assign _0155_ = pk_rsp_wr_cnt == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6245" *) 2'b10;
  assign is_last_loop = rd_loop_cnt_inc >= (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1402" *) rd_loop_cnt_limit;
  assign is_base_wrap = pk_rsp_wr_base_inc[12:8] >= (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7319" *) pixel_bank;
  assign is_addr_wrap = pk_rsp_wr_addr_inc[13:8] >= (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7978" *) pixel_bank;
  assign data_planar0_p0_cur_flag[0] = data_planar0_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2613" *) pad_left_d1;
  assign data_planar0_p0_cur_flag[1] = data_planar0_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2614" *) data_width_mark_1;
  assign data_planar0_p0_cur_flag[2] = data_planar0_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2615" *) data_width_mark_2;
  assign data_planar0_p1_cur_flag[0] = data_planar0_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2623" *) pad_left_d1;
  assign data_planar0_p1_cur_flag[1] = data_planar0_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2624" *) data_width_mark_1;
  assign data_planar0_p1_cur_flag[2] = data_planar0_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2625" *) data_width_mark_2;
  assign data_planar1_p0_cur_flag[0] = data_planar1_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2633" *) pad_left_d1;
  assign data_planar1_p0_cur_flag[1] = data_planar1_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2634" *) data_width_mark_1;
  assign data_planar1_p0_cur_flag[2] = data_planar1_p0_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2635" *) data_width_mark_2;
  assign data_planar1_p1_cur_flag[0] = data_planar1_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2643" *) pad_left_d1;
  assign data_planar1_p1_cur_flag[1] = data_planar1_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2644" *) data_width_mark_1;
  assign data_planar1_p1_cur_flag[2] = data_planar1_p1_cnt_w > (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2645" *) data_width_mark_2;
  assign is_1st_height = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1259" *) _0373_;
  assign _0157_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1574" *) rd_planar_cnt;
  assign _0158_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1580" *) pixel_planar;
  assign _0159_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1650" *) rd_pburst_cnt;
  assign _0160_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *) is_last_loop;
  assign _0161_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *) img_pd[0];
  assign _0162_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *) data_planar0_p1_flag[0];
  assign _0163_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *) _0376_;
  assign _0164_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *) data_planar0_p1_flag[1];
  assign _0165_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2715" *) data_planar0_p0_zero_mask;
  assign _0166_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2725" *) data_planar0_p0_cur_flag[0];
  assign _0167_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2728" *) data_planar0_p0_cur_flag[1];
  assign _0168_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2733" *) data_planar0_p1_zero_mask;
  assign _0169_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *) data_planar1_p1_flag[0];
  assign _0170_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *) _0379_;
  assign _0171_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *) data_planar1_p1_flag[1];
  assign _0172_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2749" *) data_planar1_p0_zero_mask;
  assign _0173_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2759" *) data_planar1_p0_cur_flag[0];
  assign _0174_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2762" *) data_planar1_p0_cur_flag[1];
  assign _0175_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2767" *) data_planar1_p1_zero_mask;
  assign _0176_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:484" *) is_running_d1;
  assign _0177_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5097" *) pk_rsp_early_end;
  assign _0178_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5499" *) rd_planar_d3;
  assign _0179_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5565" *) pixel_packed_10b;
  assign _0180_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) pk_rsp_wr_w_offset[1];
  assign _0181_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) pixel_data_expand;
  assign _0182_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *) _0375_;
  assign _0183_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7693" *) pk_rsp_cur_sub_h_end;
  assign _0184_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1409" *) is_last_loop;
  assign _0185_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1573" *) is_last_planar;
  assign is_last_planar = _0158_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1580" *) rd_planar_cnt;
  assign _0186_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1649" *) is_last_pburst;
  assign _0187_ = _0160_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1657" *) _0161_;
  assign rd_vld = sg2pack_img_pvld | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1732" *) rd_local_vld;
  assign rd_pburst_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1800" *) rd_vld;
  assign rd_planar_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1807" *) _0094_;
  assign rd_loop_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1813" *) rd_planar_end;
  assign rd_height_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1819" *) rd_line_end;
  assign rd_planar0_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1953" *) _0102_;
  assign rd_planar1_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1954" *) _0103_;
  assign _0188_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2655" *) rd_planar0_line_end;
  assign _0189_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2667" *) rd_planar1_line_end;
  assign _0190_ = data_planar0_p0_lp_mask | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2715" *) data_planar0_p0_rp_mask;
  assign _0191_ = data_planar0_p1_lp_mask | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2733" *) data_planar0_p1_rp_mask;
  assign _0192_ = data_planar1_p0_lp_mask | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2749" *) data_planar1_p0_rp_mask;
  assign _0193_ = data_planar1_p1_lp_mask | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2767" *) data_planar1_p1_rp_mask;
  assign pk_rsp_pipe_sel = _0158_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5480" *) _0117_;
  assign _0194_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5499" *) _0178_;
  assign _0195_ = pixel_data_shrink | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5566" *) _0121_;
  assign _0196_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6061" *) rd_p0_zero_mask_d3[0];
  assign _0197_ = _0196_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6061" *) rd_p0_pad_mask_d3[0];
  assign _0198_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6063" *) rd_p0_zero_mask_d3[4];
  assign _0199_ = _0198_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6063" *) rd_p0_pad_mask_d3[4];
  assign _0200_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6065" *) rd_p0_zero_mask_d3[8];
  assign _0201_ = _0200_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6065" *) rd_p0_pad_mask_d3[8];
  assign _0202_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6067" *) rd_p0_zero_mask_d3[12];
  assign _0203_ = _0202_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6067" *) rd_p0_pad_mask_d3[12];
  assign _0204_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6069" *) rd_p0_zero_mask_d3[16];
  assign _0205_ = _0204_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6069" *) rd_p0_pad_mask_d3[16];
  assign _0206_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6071" *) rd_p0_zero_mask_d3[20];
  assign _0207_ = _0206_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6071" *) rd_p0_pad_mask_d3[20];
  assign _0208_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6073" *) rd_p0_zero_mask_d3[24];
  assign _0209_ = _0208_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6073" *) rd_p0_pad_mask_d3[24];
  assign _0210_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6075" *) rd_p0_zero_mask_d3[28];
  assign _0211_ = _0210_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6075" *) rd_p0_pad_mask_d3[28];
  assign _0212_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6077" *) rd_p1_zero_mask_d3[0];
  assign _0213_ = _0212_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6077" *) rd_p1_pad_mask_d3[0];
  assign _0214_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6079" *) rd_p1_zero_mask_d3[4];
  assign _0215_ = _0214_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6079" *) rd_p1_pad_mask_d3[4];
  assign _0216_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6081" *) rd_p1_zero_mask_d3[8];
  assign _0217_ = _0216_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6081" *) rd_p1_pad_mask_d3[8];
  assign _0218_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6083" *) rd_p1_zero_mask_d3[12];
  assign _0219_ = _0218_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6083" *) rd_p1_pad_mask_d3[12];
  assign _0220_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6085" *) rd_p1_zero_mask_d3[16];
  assign _0221_ = _0220_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6085" *) rd_p1_pad_mask_d3[16];
  assign _0222_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6087" *) rd_p1_zero_mask_d3[20];
  assign _0223_ = _0222_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6087" *) rd_p1_pad_mask_d3[20];
  assign _0224_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6089" *) rd_p1_zero_mask_d3[24];
  assign _0225_ = _0224_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6089" *) rd_p1_pad_mask_d3[24];
  assign _0226_ = _0179_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6091" *) rd_p1_zero_mask_d3[28];
  assign _0227_ = _0226_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6091" *) rd_p1_pad_mask_d3[28];
  assign _0228_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6100" *) rd_p0_zero_mask_d3[0];
  assign _0229_ = _0228_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6100" *) rd_p0_pad_mask_d3[0];
  assign _0230_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6102" *) rd_p0_zero_mask_d3[1];
  assign _0231_ = _0230_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6102" *) rd_p0_pad_mask_d3[1];
  assign _0232_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6104" *) rd_p0_zero_mask_d3[2];
  assign _0233_ = _0232_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6104" *) rd_p0_pad_mask_d3[2];
  assign _0234_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6106" *) rd_p0_zero_mask_d3[3];
  assign _0235_ = _0234_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6106" *) rd_p0_pad_mask_d3[3];
  assign _0236_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6108" *) rd_p0_zero_mask_d3[4];
  assign _0237_ = _0236_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6108" *) rd_p0_pad_mask_d3[4];
  assign _0238_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6110" *) rd_p0_zero_mask_d3[5];
  assign _0239_ = _0238_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6110" *) rd_p0_pad_mask_d3[5];
  assign _0240_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6112" *) rd_p0_zero_mask_d3[6];
  assign _0241_ = _0240_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6112" *) rd_p0_pad_mask_d3[6];
  assign _0242_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6114" *) rd_p0_zero_mask_d3[7];
  assign _0243_ = _0242_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6114" *) rd_p0_pad_mask_d3[7];
  assign _0244_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6116" *) rd_p0_zero_mask_d3[8];
  assign _0245_ = _0244_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6116" *) rd_p0_pad_mask_d3[8];
  assign _0246_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6118" *) rd_p0_zero_mask_d3[9];
  assign _0247_ = _0246_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6118" *) rd_p0_pad_mask_d3[9];
  assign _0248_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6120" *) rd_p0_zero_mask_d3[10];
  assign _0249_ = _0248_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6120" *) rd_p0_pad_mask_d3[10];
  assign _0250_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6122" *) rd_p0_zero_mask_d3[11];
  assign _0251_ = _0250_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6122" *) rd_p0_pad_mask_d3[11];
  assign _0252_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6124" *) rd_p0_zero_mask_d3[12];
  assign _0253_ = _0252_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6124" *) rd_p0_pad_mask_d3[12];
  assign _0254_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6126" *) rd_p0_zero_mask_d3[13];
  assign _0255_ = _0254_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6126" *) rd_p0_pad_mask_d3[13];
  assign _0256_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6128" *) rd_p0_zero_mask_d3[14];
  assign _0257_ = _0256_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6128" *) rd_p0_pad_mask_d3[14];
  assign _0258_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6130" *) rd_p0_zero_mask_d3[15];
  assign _0259_ = _0258_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6130" *) rd_p0_pad_mask_d3[15];
  assign _0260_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6132" *) rd_p0_zero_mask_d3[16];
  assign _0261_ = _0260_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6132" *) rd_p0_pad_mask_d3[16];
  assign _0262_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6134" *) rd_p0_zero_mask_d3[17];
  assign _0263_ = _0262_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6134" *) rd_p0_pad_mask_d3[17];
  assign _0264_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6136" *) rd_p0_zero_mask_d3[18];
  assign _0265_ = _0264_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6136" *) rd_p0_pad_mask_d3[18];
  assign _0266_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6138" *) rd_p0_zero_mask_d3[19];
  assign _0267_ = _0266_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6138" *) rd_p0_pad_mask_d3[19];
  assign _0268_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6140" *) rd_p0_zero_mask_d3[20];
  assign _0269_ = _0268_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6140" *) rd_p0_pad_mask_d3[20];
  assign _0270_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6142" *) rd_p0_zero_mask_d3[21];
  assign _0271_ = _0270_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6142" *) rd_p0_pad_mask_d3[21];
  assign _0272_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6144" *) rd_p0_zero_mask_d3[22];
  assign _0273_ = _0272_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6144" *) rd_p0_pad_mask_d3[22];
  assign _0274_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6146" *) rd_p0_zero_mask_d3[23];
  assign _0275_ = _0274_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6146" *) rd_p0_pad_mask_d3[23];
  assign _0276_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6148" *) rd_p0_zero_mask_d3[24];
  assign _0277_ = _0276_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6148" *) rd_p0_pad_mask_d3[24];
  assign _0278_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6150" *) rd_p0_zero_mask_d3[25];
  assign _0279_ = _0278_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6150" *) rd_p0_pad_mask_d3[25];
  assign _0280_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6152" *) rd_p0_zero_mask_d3[26];
  assign _0281_ = _0280_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6152" *) rd_p0_pad_mask_d3[26];
  assign _0282_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6154" *) rd_p0_zero_mask_d3[27];
  assign _0283_ = _0282_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6154" *) rd_p0_pad_mask_d3[27];
  assign _0284_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6156" *) rd_p0_zero_mask_d3[28];
  assign _0285_ = _0284_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6156" *) rd_p0_pad_mask_d3[28];
  assign _0286_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6158" *) rd_p0_zero_mask_d3[29];
  assign _0287_ = _0286_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6158" *) rd_p0_pad_mask_d3[29];
  assign _0288_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6160" *) rd_p0_zero_mask_d3[30];
  assign _0289_ = _0288_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6160" *) rd_p0_pad_mask_d3[30];
  assign _0290_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6162" *) rd_p0_zero_mask_d3[31];
  assign _0291_ = _0290_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6162" *) rd_p0_pad_mask_d3[31];
  assign _0292_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6164" *) rd_p1_zero_mask_d3[0];
  assign _0293_ = _0292_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6164" *) rd_p1_pad_mask_d3[0];
  assign _0294_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6166" *) rd_p1_zero_mask_d3[1];
  assign _0295_ = _0294_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6166" *) rd_p1_pad_mask_d3[1];
  assign _0296_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6168" *) rd_p1_zero_mask_d3[2];
  assign _0297_ = _0296_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6168" *) rd_p1_pad_mask_d3[2];
  assign _0298_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6170" *) rd_p1_zero_mask_d3[3];
  assign _0299_ = _0298_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6170" *) rd_p1_pad_mask_d3[3];
  assign _0300_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6172" *) rd_p1_zero_mask_d3[4];
  assign _0301_ = _0300_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6172" *) rd_p1_pad_mask_d3[4];
  assign _0302_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6174" *) rd_p1_zero_mask_d3[5];
  assign _0303_ = _0302_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6174" *) rd_p1_pad_mask_d3[5];
  assign _0304_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6176" *) rd_p1_zero_mask_d3[6];
  assign _0305_ = _0304_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6176" *) rd_p1_pad_mask_d3[6];
  assign _0306_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6178" *) rd_p1_zero_mask_d3[7];
  assign _0307_ = _0306_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6178" *) rd_p1_pad_mask_d3[7];
  assign _0308_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6180" *) rd_p1_zero_mask_d3[8];
  assign _0309_ = _0308_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6180" *) rd_p1_pad_mask_d3[8];
  assign _0310_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6182" *) rd_p1_zero_mask_d3[9];
  assign _0311_ = _0310_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6182" *) rd_p1_pad_mask_d3[9];
  assign _0312_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6184" *) rd_p1_zero_mask_d3[10];
  assign _0313_ = _0312_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6184" *) rd_p1_pad_mask_d3[10];
  assign _0314_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6186" *) rd_p1_zero_mask_d3[11];
  assign _0315_ = _0314_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6186" *) rd_p1_pad_mask_d3[11];
  assign _0316_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6188" *) rd_p1_zero_mask_d3[12];
  assign _0317_ = _0316_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6188" *) rd_p1_pad_mask_d3[12];
  assign _0318_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6190" *) rd_p1_zero_mask_d3[13];
  assign _0319_ = _0318_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6190" *) rd_p1_pad_mask_d3[13];
  assign _0320_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6192" *) rd_p1_zero_mask_d3[14];
  assign _0321_ = _0320_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6192" *) rd_p1_pad_mask_d3[14];
  assign _0322_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6194" *) rd_p1_zero_mask_d3[15];
  assign _0323_ = _0322_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6194" *) rd_p1_pad_mask_d3[15];
  assign _0324_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6196" *) rd_p1_zero_mask_d3[16];
  assign _0325_ = _0324_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6196" *) rd_p1_pad_mask_d3[16];
  assign _0326_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6198" *) rd_p1_zero_mask_d3[17];
  assign _0327_ = _0326_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6198" *) rd_p1_pad_mask_d3[17];
  assign _0328_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6200" *) rd_p1_zero_mask_d3[18];
  assign _0329_ = _0328_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6200" *) rd_p1_pad_mask_d3[18];
  assign _0330_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6202" *) rd_p1_zero_mask_d3[19];
  assign _0331_ = _0330_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6202" *) rd_p1_pad_mask_d3[19];
  assign _0332_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6204" *) rd_p1_zero_mask_d3[20];
  assign _0333_ = _0332_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6204" *) rd_p1_pad_mask_d3[20];
  assign _0334_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6206" *) rd_p1_zero_mask_d3[21];
  assign _0335_ = _0334_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6206" *) rd_p1_pad_mask_d3[21];
  assign _0336_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6208" *) rd_p1_zero_mask_d3[22];
  assign _0337_ = _0336_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6208" *) rd_p1_pad_mask_d3[22];
  assign _0338_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6210" *) rd_p1_zero_mask_d3[23];
  assign _0339_ = _0338_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6210" *) rd_p1_pad_mask_d3[23];
  assign _0340_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6212" *) rd_p1_zero_mask_d3[24];
  assign _0341_ = _0340_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6212" *) rd_p1_pad_mask_d3[24];
  assign _0342_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6214" *) rd_p1_zero_mask_d3[25];
  assign _0343_ = _0342_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6214" *) rd_p1_pad_mask_d3[25];
  assign _0344_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6216" *) rd_p1_zero_mask_d3[26];
  assign _0345_ = _0344_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6216" *) rd_p1_pad_mask_d3[26];
  assign _0346_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6218" *) rd_p1_zero_mask_d3[27];
  assign _0347_ = _0346_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6218" *) rd_p1_pad_mask_d3[27];
  assign _0348_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6220" *) rd_p1_zero_mask_d3[28];
  assign _0349_ = _0348_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6220" *) rd_p1_pad_mask_d3[28];
  assign _0350_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6222" *) rd_p1_zero_mask_d3[29];
  assign _0351_ = _0350_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6222" *) rd_p1_pad_mask_d3[29];
  assign _0352_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6224" *) rd_p1_zero_mask_d3[30];
  assign _0353_ = _0352_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6224" *) rd_p1_pad_mask_d3[30];
  assign _0354_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6226" *) rd_p1_zero_mask_d3[31];
  assign _0355_ = _0354_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6226" *) rd_p1_pad_mask_d3[31];
  assign _0356_ = _0122_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6259" *) _0123_;
  assign _0357_ = _0356_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6260" *) _0124_;
  assign _0358_ = _0357_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6261" *) _0125_;
  assign pk_rsp_data_h0 = _0358_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6262" *) _0126_;
  assign _0359_ = _0127_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6286" *) _0128_;
  assign _0360_ = _0359_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6287" *) _0129_;
  assign _0361_ = _0360_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6288" *) _0130_;
  assign pk_rsp_pad_mask_h0 = _0361_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6289" *) _0131_;
  assign _0156_ = pk_rsp_data_h1_en | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6686" *) is_first_running;
  assign _0362_ = pixel_packed_10b | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *) _0182_;
  assign _0363_ = _0133_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7051" *) _0134_;
  assign _0364_ = _0363_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7052" *) _0135_;
  assign pk_rsp_mn_data_h1 = _0364_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7053" *) _0136_;
  assign _0365_ = _0137_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7063" *) _0138_;
  assign _0366_ = _0365_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7064" *) _0139_;
  assign _0367_ = _0366_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7065" *) _0140_;
  assign _0368_ = _0367_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7066" *) _0141_;
  assign _0369_ = _0368_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7067" *) _0142_;
  assign _0370_ = _0369_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7068" *) _0143_;
  assign pk_rsp_mn_data_h0 = _0370_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7069" *) _0144_;
  assign pk_rsp_wr_base_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7342" *) pk_rsp_data_updt;
  assign _0371_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7507" *) pk_rsp_cur_sub_h_end;
  assign pk_rsp_wr_h_offset_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7515" *) _0146_;
  assign _0372_ = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7692" *) _0147_;
  assign pk_rsp_wr_w_offset_en = is_first_running | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7700" *) pk_rsp_wr_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pack_is_done <= 1'b1;
    else
      pack_is_done <= pack_is_done_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_data_slices <= 4'b0000;
    else
      pk_out_data_slices <= _0019_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_data_entries <= 12'b000000000000;
    else
      pk_out_data_entries <= _0016_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_data_updt <= 1'b0;
    else
      pk_out_data_updt <= pk_rsp_data_updt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_hsel <= 1'b0;
    else
      pk_out_hsel <= _0022_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_addr <= 12'b000000000000;
    else
      pk_out_addr <= _0015_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_wr_w_offset_ori <= 14'b00000000000000;
    else
      pk_rsp_wr_w_offset_ori <= _0040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_wr_w_offset <= 14'b00000000000000;
    else
      pk_rsp_wr_w_offset <= _0039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_wr_h_offset <= 12'b000000000000;
    else
      pk_rsp_wr_h_offset <= _0038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_wr_base <= 12'b000000000000;
    else
      pk_rsp_wr_base <= _0036_;
  always @(posedge nvdla_core_clk)
      pk_mn_out_data_h0 <= _0013_;
  always @(posedge nvdla_core_clk)
      pk_mn_out_data_h1 <= _0014_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mn_mask_uv_lo_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mn_mask_uv_lo_d1 <= mn_mask_uv_lo;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mn_mask_y_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mn_mask_y_d1 <= _0011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_pad_mask_h0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      pk_out_pad_mask_h0 <= _0025_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_pad_mask_h1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      pk_out_pad_mask_h1 <= _0026_;
  always @(posedge nvdla_core_clk)
      pk_out_data_h0 <= _0017_;
  always @(posedge nvdla_core_clk)
      pk_out_data_h1 <= _0018_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mask_pad_planar1_c1_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mask_pad_planar1_c1_d1 <= pad_mask_l1_hi;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mask_pad_planar1_c0_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mask_pad_planar1_c0_d1 <= pad_mask_l1_lo;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mask_pad_planar0_c0_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mask_pad_planar0_c0_d1 <= _0010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_planar1_c1_d1 <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      pk_rsp_planar1_c1_d1 <= dat_l1_hi;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_planar1_c0_d1 <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      pk_rsp_planar1_c0_d1 <= dat_l1_lo;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_planar0_c0_d1 <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      pk_rsp_planar0_c0_d1 <= _0033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_ext128 <= 1'b0;
    else
      pk_out_ext128 <= _0020_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_ext64 <= 1'b0;
    else
      pk_out_ext64 <= _0021_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_uint <= 1'b0;
    else
      pk_out_uint <= _0028_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_mean <= 1'b0;
    else
      pk_out_mean <= _0024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_mask <= 4'b0000;
    else
      pk_out_mask <= _0023_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_sub_h <= 3'b000;
    else
      pk_out_sub_h <= _0027_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_out_vld <= 1'b0;
    else
      pk_out_vld <= pk_rsp_wr_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_wr_cnt <= 2'b00;
    else
      pk_rsp_wr_cnt <= _0037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_layer_end_d1 <= 1'b0;
    else
      pk_rsp_layer_end_d1 <= _0030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_1st_height_d1 <= 1'b0;
    else
      pk_rsp_1st_height_d1 <= _0029_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_one_line_end_d1 <= 1'b0;
    else
      pk_rsp_one_line_end_d1 <= _0032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_loop_end_d1 <= 1'b0;
    else
      pk_rsp_loop_end_d1 <= _0031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_sub_h_end_d1 <= 1'b0;
    else
      pk_rsp_sub_h_end_d1 <= _0035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_sub_h_d1 <= 3'b000;
    else
      pk_rsp_sub_h_d1 <= _0034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pk_rsp_vld_d1 <= 1'b0;
    else
      pk_rsp_vld_d1 <= pk_rsp_vld_d1_w;
  always @(posedge nvdla_core_clk)
      rd_p1_zero_mask_d3 <= _0072_;
  always @(posedge nvdla_core_clk)
      rd_p0_zero_mask_d3 <= _0063_;
  always @(posedge nvdla_core_clk)
      rd_p1_pad_mask_d3 <= _0067_;
  always @(posedge nvdla_core_clk)
      rd_p0_pad_mask_d3 <= _0058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_layer_end_d3 <= 1'b0;
    else
      rd_layer_end_d3 <= _0047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_1st_height_d3 <= 1'b0;
    else
      rd_1st_height_d3 <= _0043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_one_line_end_d3 <= 1'b0;
    else
      rd_one_line_end_d3 <= _0054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_loop_end_d3 <= 1'b0;
    else
      rd_loop_end_d3 <= _0051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_end_d3 <= 1'b0;
    else
      rd_sub_h_end_d3 <= _0083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_d3 <= 3'b000;
    else
      rd_sub_h_d3 <= _0080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_planar_d3 <= 1'b0;
    else
      rd_planar_d3 <= _0077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_vld_d3 <= 1'b0;
    else
      rd_vld_d3 <= rd_vld_d2;
  always @(posedge nvdla_core_clk)
      rd_p1_zero_mask_d2 <= _0071_;
  always @(posedge nvdla_core_clk)
      rd_p0_zero_mask_d2 <= _0062_;
  always @(posedge nvdla_core_clk)
      rd_p1_pad_mask_d2 <= _0066_;
  always @(posedge nvdla_core_clk)
      rd_p0_pad_mask_d2 <= _0057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_layer_end_d2 <= 1'b0;
    else
      rd_layer_end_d2 <= _0046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_1st_height_d2 <= 1'b0;
    else
      rd_1st_height_d2 <= _0042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_one_line_end_d2 <= 1'b0;
    else
      rd_one_line_end_d2 <= _0053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_loop_end_d2 <= 1'b0;
    else
      rd_loop_end_d2 <= _0050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_end_d2 <= 1'b0;
    else
      rd_sub_h_end_d2 <= _0082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_d2 <= 3'b000;
    else
      rd_sub_h_d2 <= _0079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_planar_d2 <= 1'b0;
    else
      rd_planar_d2 <= _0076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_vld_d2 <= 1'b0;
    else
      rd_vld_d2 <= rd_vld_d1;
  always @(posedge nvdla_core_clk)
      rd_p1_zero_mask_d1 <= _0070_;
  always @(posedge nvdla_core_clk)
      rd_p0_zero_mask_d1 <= _0061_;
  always @(posedge nvdla_core_clk)
      rd_p1_pad_mask_d1 <= _0065_;
  always @(posedge nvdla_core_clk)
      rd_p0_pad_mask_d1 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_layer_end_d1 <= 1'b0;
    else
      rd_layer_end_d1 <= _0045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_1st_height_d1 <= 1'b0;
    else
      rd_1st_height_d1 <= _0041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_one_line_end_d1 <= 1'b0;
    else
      rd_one_line_end_d1 <= _0052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_loop_end_d1 <= 1'b0;
    else
      rd_loop_end_d1 <= _0049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_end_d1 <= 1'b0;
    else
      rd_sub_h_end_d1 <= _0081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_h_d1 <= 3'b000;
    else
      rd_sub_h_d1 <= _0078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_planar_d1 <= 1'b0;
    else
      rd_planar_d1 <= _0075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar1_p1_flag <= 3'b000;
    else
      data_planar1_p1_flag <= _0005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar0_p1_flag <= 3'b000;
    else
      data_planar0_p1_flag <= _0002_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar1_cur_cnt <= 14'b00000000000000;
    else
      data_planar1_cur_cnt <= _0004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar0_cur_cnt <= 14'b00000000000000;
    else
      data_planar0_cur_cnt <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p1_addr_d1 <= 8'b00000000;
    else
      rd_p1_addr_d1 <= _0064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p0_addr_d1 <= 8'b00000000;
    else
      rd_p0_addr_d1 <= _0055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p1_planar1_idx <= 7'b0000000;
    else
      rd_p1_planar1_idx <= _0069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p1_planar0_idx <= 7'b0000000;
    else
      rd_p1_planar0_idx <= _0068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p0_planar1_idx <= 7'b0000000;
    else
      rd_p0_planar1_idx <= _0060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p0_planar0_idx <= 7'b0000000;
    else
      rd_p0_planar0_idx <= _0059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p1_vld_d1 <= 1'b0;
    else
      rd_p1_vld_d1 <= rd_p1_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_p0_vld_d1 <= 1'b0;
    else
      rd_p0_vld_d1 <= rd_p0_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_vld_d1 <= 1'b0;
    else
      rd_vld_d1 <= rd_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_local_vld <= 1'b0;
    else
      rd_local_vld <= rd_local_vld_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pburst_cnt <= 1'b0;
    else
      rd_pburst_cnt <= _0073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_planar_cnt <= 1'b0;
    else
      rd_planar_cnt <= _0074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_loop_cnt <= 3'b000;
    else
      rd_loop_cnt <= _0048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_height_cnt <= 13'b0000000000000;
    else
      rd_height_cnt <= _0044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar1_add <= 6'b000000;
    else
      data_planar1_add <= _0003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_planar0_add <= 6'b000000;
    else
      data_planar0_add <= _0000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      zero_planar1_mask_sft <= 5'b00000;
    else
      zero_planar1_mask_sft <= _0087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      zero_planar0_mask_sft <= 5'b00000;
    else
      zero_planar0_mask_sft <= _0086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rp_planar1_mask_sft <= 5'b00000;
    else
      rp_planar1_mask_sft <= _0085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rp_planar0_mask_sft <= 5'b00000;
    else
      rp_planar0_mask_sft <= _0084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lp_planar1_mask_sft <= 5'b00000;
    else
      lp_planar1_mask_sft <= _0009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lp_planar0_mask_sft <= 5'b00000;
    else
      lp_planar0_mask_sft <= _0008_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_width_mark_2 <= 14'b00000000000000;
    else
      data_width_mark_2 <= _0007_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_width_mark_1 <= 14'b00000000000000;
    else
      data_width_mark_1 <= _0006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pad_left_d1 <= 5'b00000;
    else
      pad_left_d1 <= _0012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      is_running_d1 <= 1'b0;
    else
      is_running_d1 <= is_running;
  assign _0019_ = pk_rsp_data_updt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8343" *) pk_rsp_data_slices : pk_out_data_slices;
  assign _0016_ = pk_rsp_data_updt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8282" *) pk_rsp_data_entries : pk_out_data_entries;
  assign _0022_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8061" *) pk_rsp_wr_w_offset[1] : pk_out_hsel;
  assign _0015_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8000" *) pk_rsp_wr_addr : pk_out_addr;
  assign _0040_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7768" *) pk_rsp_wr_w_offset_w : pk_rsp_wr_w_offset_ori;
  assign _0039_ = pk_rsp_wr_w_offset_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7707" *) pk_rsp_wr_w_offset_w : pk_rsp_wr_w_offset;
  assign _0038_ = pk_rsp_wr_h_offset_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7521" *) pk_rsp_wr_h_offset_w : pk_rsp_wr_h_offset;
  assign _0036_ = pk_rsp_wr_base_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7348" *) pk_rsp_wr_base_w : pk_rsp_wr_base;
  assign _0013_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7270" *) pk_rsp_mn_data_h0 : pk_mn_out_data_h0;
  assign _0014_ = pk_rsp_mn_data_h1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7260" *) pk_rsp_mn_data_h1 : pk_mn_out_data_h1;
  assign mn_mask_uv_lo = mn_mask_uv_0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7141" *) { rd_p1_zero_mask_d3, rd_p0_zero_mask_d3 } : mn_mask_uv_lo_d1;
  assign _0011_ = mn_mask_y_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7080" *) { rd_p1_zero_mask_d3, rd_p0_zero_mask_d3 } : mn_mask_y_d1;
  assign _0025_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6747" *) pk_rsp_pad_mask_h0 : pk_out_pad_mask_h0;
  assign _0026_ = _0156_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6686" *) pk_rsp_pad_mask_h1 : pk_out_pad_mask_h1;
  assign _0017_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6673" *) pk_rsp_data_h0 : pk_out_data_h0;
  assign _0018_ = pk_rsp_data_h1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6663" *) pk_rsp_data_h1 : pk_out_data_h1;
  assign pad_mask_l1_hi = pk_rsp_planar1_c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6605" *) { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 } : mask_pad_planar1_c1_d1;
  assign pad_mask_l1_lo = mn_mask_uv_0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6544" *) { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 } : mask_pad_planar1_c0_d1;
  assign _0010_ = mn_mask_y_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6483" *) { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 } : mask_pad_planar0_c0_d1;
  assign dat_l1_hi = pk_rsp_planar1_c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6422" *) pk_rsp_dat_mnorm : pk_rsp_planar1_c1_d1;
  assign dat_l1_lo = mn_mask_uv_0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6361" *) pk_rsp_dat_mnorm : pk_rsp_planar1_c0_d1;
  assign _0033_ = mn_mask_y_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6300" *) pk_rsp_dat_mnorm : pk_rsp_planar0_c0_d1;
  assign _0020_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5884" *) pk_rsp_wr_ext128 : pk_out_ext128;
  assign _0021_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5823" *) pk_rsp_wr_ext64 : pk_out_ext64;
  assign _0028_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5762" *) pixel_uint : pk_out_uint;
  assign _0024_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5701" *) sg2pack_mn_enable : pk_out_mean;
  assign _0023_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5640" *) pk_rsp_wr_mask : pk_out_mask;
  assign _0027_ = pk_rsp_wr_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5579" *) pk_rsp_cur_sub_h : pk_out_sub_h;
  assign _0037_ = rd_vld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5506" *) pk_rsp_wr_cnt_w : pk_rsp_wr_cnt;
  assign _0030_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5414" *) rd_layer_end_d3 : pk_rsp_layer_end_d1;
  assign _0029_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5353" *) rd_1st_height_d3 : pk_rsp_1st_height_d1;
  assign _0032_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5292" *) rd_one_line_end_d3 : pk_rsp_one_line_end_d1;
  assign _0031_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5231" *) rd_loop_end_d3 : pk_rsp_loop_end_d1;
  assign _0035_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5170" *) rd_sub_h_end_d3 : pk_rsp_sub_h_end_d1;
  assign _0034_ = pk_rsp_vld_d1_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5109" *) rd_sub_h_d3 : pk_rsp_sub_h_d1;
  assign _0072_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5075" *) rd_p1_zero_mask_d2 : rd_p1_zero_mask_d3;
  assign _0063_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5065" *) rd_p0_zero_mask_d2 : rd_p0_zero_mask_d3;
  assign _0067_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5055" *) rd_p1_pad_mask_d2 : rd_p1_pad_mask_d3;
  assign _0058_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5045" *) rd_p0_pad_mask_d2 : rd_p0_pad_mask_d3;
  assign _0047_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4987" *) rd_layer_end_d2 : rd_layer_end_d3;
  assign _0043_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4926" *) rd_1st_height_d2 : rd_1st_height_d3;
  assign _0054_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4865" *) rd_one_line_end_d2 : rd_one_line_end_d3;
  assign _0051_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4804" *) rd_loop_end_d2 : rd_loop_end_d3;
  assign _0083_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4743" *) rd_sub_h_end_d2 : rd_sub_h_end_d3;
  assign _0080_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4682" *) rd_sub_h_d2 : rd_sub_h_d3;
  assign _0077_ = rd_vld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4621" *) rd_planar_d2 : rd_planar_d3;
  assign _0071_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4601" *) rd_p1_zero_mask_d1 : rd_p1_zero_mask_d2;
  assign _0062_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4591" *) rd_p0_zero_mask_d1 : rd_p0_zero_mask_d2;
  assign _0066_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4581" *) rd_p1_pad_mask_d1 : rd_p1_pad_mask_d2;
  assign _0057_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4571" *) rd_p0_pad_mask_d1 : rd_p0_pad_mask_d2;
  assign _0046_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4513" *) rd_layer_end_d1 : rd_layer_end_d2;
  assign _0042_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4452" *) rd_1st_height_d1 : rd_1st_height_d2;
  assign _0053_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4391" *) rd_one_line_end_d1 : rd_one_line_end_d2;
  assign _0050_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4330" *) rd_loop_end_d1 : rd_loop_end_d2;
  assign _0082_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4269" *) rd_sub_h_end_d1 : rd_sub_h_end_d2;
  assign _0079_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4208" *) rd_sub_h_d1 : rd_sub_h_d2;
  assign _0076_ = rd_vld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:4147" *) rd_planar_d1 : rd_planar_d2;
  assign _0070_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3741" *) rd_p1_zero_mask : rd_p1_zero_mask_d1;
  assign _0061_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3731" *) rd_p0_zero_mask : rd_p0_zero_mask_d1;
  assign _0065_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3721" *) rd_p1_pad_mask : rd_p1_pad_mask_d1;
  assign _0056_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3711" *) rd_p0_pad_mask : rd_p0_pad_mask_d1;
  assign _0045_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3653" *) _0115_ : rd_layer_end_d1;
  assign _0041_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3592" *) is_1st_height : rd_1st_height_d1;
  assign _0052_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3531" *) _0114_ : rd_one_line_end_d1;
  assign _0049_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3470" *) rd_loop_end : rd_loop_end_d1;
  assign _0081_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3409" *) rd_loop_end : rd_sub_h_end_d1;
  assign _0078_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3348" *) 3'b000 : rd_sub_h_d1;
  assign _0075_ = rd_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3287" *) rd_planar_cnt : rd_planar_d1;
  assign _0005_ = rd_planar1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3104" *) data_planar1_p1_flag_w : data_planar1_p1_flag;
  assign _0002_ = rd_planar0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:3043" *) data_planar0_p1_flag_w : data_planar0_p1_flag;
  assign _0004_ = rd_planar1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2860" *) data_planar1_cur_cnt_w : data_planar1_cur_cnt;
  assign _0001_ = rd_planar0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2799" *) data_planar0_cur_cnt_w : data_planar0_cur_cnt;
  assign _0064_ = rd_p1_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2531" *) rd_p1_addr : rd_p1_addr_d1;
  assign _0055_ = rd_p0_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2470" *) rd_p0_addr : rd_p0_addr_d1;
  assign _0069_ = rd_planar1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2165" *) rd_p1_planar1_idx_w : rd_p1_planar1_idx;
  assign _0068_ = rd_planar0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2104" *) rd_p1_planar0_idx_w : rd_p1_planar0_idx;
  assign _0060_ = rd_planar1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2043" *) rd_p0_planar1_idx_w : rd_p0_planar1_idx;
  assign _0059_ = rd_planar0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1982" *) rd_p0_planar0_idx_w : rd_p0_planar0_idx;
  assign _0073_ = rd_pburst_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1669" *) rd_pburst_cnt_w : rd_pburst_cnt;
  assign _0074_ = rd_planar_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1586" *) rd_planar_cnt_w : rd_planar_cnt;
  assign _0048_ = rd_loop_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1416" *) rd_loop_cnt_w : rd_loop_cnt;
  assign _0044_ = rd_height_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1278" *) rd_height_cnt_w : rd_height_cnt;
  assign _0003_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1190" *) data_planar1_add_w : data_planar1_add;
  assign _0000_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1129" *) data_planar0_add_w : data_planar0_add;
  assign _0087_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1068" *) zero_planar1_mask_sft_w : zero_planar1_mask_sft;
  assign _0086_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1007" *) zero_planar0_mask_sft_w : zero_planar0_mask_sft;
  assign _0085_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:946" *) rp_planar1_mask_sft_w : rp_planar1_mask_sft;
  assign _0084_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:885" *) rp_planar0_mask_sft_w : rp_planar0_mask_sft;
  assign _0009_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:824" *) lp_planar1_mask_sft_w : lp_planar1_mask_sft;
  assign _0008_ = is_first_running ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:763" *) lp_planar0_mask_sft_w : lp_planar0_mask_sft;
  assign _0007_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:702" *) data_width_mark_2_w : data_width_mark_2;
  assign _0006_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:641" *) data_width_mark_1_w : data_width_mark_1;
  assign _0012_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:580" *) reg2dp_pad_left : pad_left_d1;
  assign _0373_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1259" *) { rd_height_cnt[0], rd_height_cnt[1], rd_height_cnt[2], rd_height_cnt[3], rd_height_cnt[4], rd_height_cnt[5], rd_height_cnt[6], rd_height_cnt[7], rd_height_cnt[8], rd_height_cnt[9], rd_height_cnt[10], rd_height_cnt[11], rd_height_cnt[12] };
  assign _0374_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6817" *) { reg2dp_datain_channel[0], reg2dp_datain_channel[1], reg2dp_datain_channel[2], reg2dp_datain_channel[3], reg2dp_datain_channel[4], reg2dp_datain_channel[5], reg2dp_datain_channel[6], reg2dp_datain_channel[7], reg2dp_datain_channel[8], reg2dp_datain_channel[9], reg2dp_datain_channel[10], reg2dp_datain_channel[11], reg2dp_datain_channel[12] };
  assign _0375_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7036" *) { pixel_precision[0], pixel_precision[1] };
  assign _0376_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2709" *) lp_planar0_mask_sft;
  assign _0377_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2712" *) rp_planar0_mask_sft;
  assign _0378_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2714" *) zero_planar0_mask_sft;
  assign _0379_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2743" *) lp_planar1_mask_sft;
  assign _0380_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2746" *) rp_planar1_mask_sft;
  assign _0381_ = 32'd4294967295 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2748" *) zero_planar1_mask_sft;
  assign data_planar0_add_w = 1'b1 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:573" *) pixel_planar0_sft;
  assign data_planar1_add_w = 1'b1 << (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:574" *) pixel_planar1_sft;
  assign lp_planar0_mask_sft_w = { pad_left_d1, 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:550" *) pixel_planar0_sft;
  assign lp_planar1_mask_sft_w = { pad_left_d1, 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:551" *) pixel_planar1_sft;
  assign rp_planar0_mask_sft_w = { data_width_mark_1[4:0], 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:558" *) pixel_planar0_sft;
  assign rp_planar1_mask_sft_w = { data_width_mark_1[4:0], 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:559" *) pixel_planar1_sft;
  assign zero_planar0_mask_sft_w = { data_width_mark_2[4:0], 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:566" *) pixel_planar0_sft;
  assign zero_planar1_mask_sft_w = { data_width_mark_2[4:0], 5'b00000 } >> (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:567" *) pixel_planar1_sft;
  assign pk_rsp_wr_base_wrap = pk_rsp_wr_base_inc[11:8] - (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7326" *) pixel_bank;
  assign pk_rsp_wr_addr_wrap = pk_rsp_wr_addr_inc[11:8] - (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7985" *) pixel_bank;
  assign rd_height_cnt_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1272" *) 13'b0000000000000 : rd_height_cnt_inc;
  assign rd_loop_cnt_w = _0184_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1410" *) 3'b000 : rd_loop_cnt_inc;
  assign rd_planar_cnt_w = _0185_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1574" *) 1'b0 : _0157_;
  assign rd_pburst_cnt_w = _0186_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1650" *) 1'b0 : _0159_;
  assign _0382_ = sg2pack_img_pvld ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1743" *) 1'b1 : rd_local_vld;
  assign _0383_ = rd_loop_end ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1743" *) 1'b0 : _0382_;
  assign rd_local_vld_w = is_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1743" *) _0383_ : 1'b0;
  assign rd_planar0_rd_mask = _0100_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1865" *) 2'b01 : 2'b11;
  assign rd_planar1_rd_mask = _0101_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1866" *) 2'b01 : 2'b11;
  assign rd_rd_mask = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1873" *) rd_planar1_rd_mask : rd_planar0_rd_mask;
  assign rd_idx_add = rd_rd_mask[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1900" *) 2'b10 : 2'b01;
  assign rd_p0_planar0_idx_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1926" *) 7'b0000000 : rd_p0_planar0_idx_inc;
  assign rd_p1_planar0_idx_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1929" *) 7'b0000001 : rd_p1_planar0_idx_inc;
  assign rd_p0_planar1_idx_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1943" *) 7'b0000000 : rd_p0_planar1_idx_inc;
  assign rd_p1_planar1_idx_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1946" *) 7'b0000001 : rd_p1_planar1_idx_inc;
  assign rd_p0_addr = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1968" *) { 1'b1, rd_p0_planar1_idx[0], rd_p0_planar1_idx[6:1] } : { 1'b0, rd_p0_planar0_idx[0], rd_p0_planar0_idx[6:1] };
  assign rd_p1_addr = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:1976" *) { 1'b1, rd_p1_planar1_idx[0], rd_p1_planar1_idx[6:1] } : { 1'b0, rd_p1_planar0_idx[0], rd_p1_planar0_idx[6:1] };
  assign data_planar0_p1_flag_w = _0188_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2657" *) 3'b000 : data_planar0_p1_cur_flag;
  assign data_planar1_p1_flag_w = _0189_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2669" *) 3'b000 : data_planar1_p1_cur_flag;
  assign _0384_ = rd_p1_vld ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2684" *) data_planar0_p1_cnt_w : data_planar0_p0_cnt_w;
  assign data_planar0_cur_cnt_w = _0188_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2684" *) 14'b00000000000000 : _0384_;
  assign _0385_ = rd_p1_vld ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2699" *) data_planar1_p1_cnt_w : data_planar1_p0_cnt_w;
  assign data_planar1_cur_cnt_w = _0189_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2699" *) 14'b00000000000000 : _0385_;
  assign _0386_ = _0104_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2710" *) _0163_ : 32'd0;
  assign data_planar0_p0_lp_mask = data_planar0_p0_cur_flag[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2710" *) _0386_ : 32'd4294967295;
  assign _0387_ = _0105_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2713" *) _0377_ : 32'd4294967295;
  assign data_planar0_p0_rp_mask = data_planar0_p0_cur_flag[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2713" *) _0387_ : 32'd0;
  assign data_planar0_p0_zero_mask = data_planar0_p0_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2714" *) _0378_ : 32'd0;
  assign _0388_ = _0106_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2726" *) _0163_ : 32'd0;
  assign data_planar0_p1_lp_mask = data_planar0_p1_cur_flag[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2726" *) _0388_ : 32'd4294967295;
  assign _0389_ = _0107_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2729" *) _0377_ : 32'd4294967295;
  assign data_planar0_p1_rp_mask = data_planar0_p1_cur_flag[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2729" *) _0389_ : 32'd0;
  assign _0390_ = data_planar0_p0_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2732" *) 32'd4294967295 : _0378_;
  assign data_planar0_p1_zero_mask = data_planar0_p1_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2732" *) _0390_ : 32'd0;
  assign _0391_ = _0108_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2744" *) _0170_ : 32'd0;
  assign data_planar1_p0_lp_mask = data_planar1_p0_cur_flag[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2744" *) _0391_ : 32'd4294967295;
  assign _0392_ = _0109_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2747" *) _0380_ : 32'd4294967295;
  assign data_planar1_p0_rp_mask = data_planar1_p0_cur_flag[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2747" *) _0392_ : 32'd0;
  assign data_planar1_p0_zero_mask = data_planar1_p0_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2748" *) _0381_ : 32'd0;
  assign _0393_ = _0110_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2760" *) _0170_ : 32'd0;
  assign data_planar1_p1_lp_mask = data_planar1_p1_cur_flag[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2760" *) _0393_ : 32'd4294967295;
  assign _0394_ = _0111_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2763" *) _0380_ : 32'd4294967295;
  assign data_planar1_p1_rp_mask = data_planar1_p1_cur_flag[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2763" *) _0394_ : 32'd0;
  assign _0395_ = data_planar1_p0_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2766" *) 32'd4294967295 : _0381_;
  assign data_planar1_p1_zero_mask = data_planar1_p1_cur_flag[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2766" *) _0395_ : 32'd0;
  assign rd_p0_pad_mask = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2780" *) data_planar1_p0_pad_mask : data_planar0_p0_pad_mask;
  assign rd_p1_pad_mask = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2781" *) data_planar1_p1_pad_mask : data_planar0_p1_pad_mask;
  assign rd_p0_zero_mask = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2782" *) data_planar1_p0_zero_mask : data_planar0_p0_zero_mask;
  assign rd_p1_zero_mask = rd_planar_cnt ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:2783" *) data_planar1_p1_zero_mask : data_planar0_p1_zero_mask;
  assign img_pd = sg2pack_img_pvld ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:474" *) sg2pack_img_pd : 11'b00000000000;
  assign pk_rsp_wr_vld = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5481" *) rd_vld_d3 : pk_rsp_vld_d1;
  assign pk_rsp_cur_sub_h = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5482" *) rd_sub_h_d3 : pk_rsp_sub_h_d1;
  assign pk_rsp_cur_sub_h_end = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5483" *) rd_sub_h_end_d3 : pk_rsp_sub_h_end_d1;
  assign pk_rsp_cur_loop_end = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5484" *) rd_loop_end_d3 : pk_rsp_loop_end_d1;
  assign pk_rsp_cur_one_line_end = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5485" *) rd_one_line_end_d3 : pk_rsp_one_line_end_d1;
  assign pk_rsp_cur_1st_height = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5486" *) rd_1st_height_d3 : pk_rsp_1st_height_d1;
  assign pk_rsp_cur_layer_end = pk_rsp_pipe_sel ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5487" *) rd_layer_end_d3 : pk_rsp_layer_end_d1;
  assign pk_rsp_wr_cnt_w = _0194_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5500" *) 2'b00 : _0089_;
  assign pk_rsp_wr_size_ori = pixel_packed_10b ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5563" *) 3'b100 : 3'b010;
  assign pk_rsp_wr_mask = pixel_packed_10b ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:5564" *) 4'b1111 : 4'b0011;
  assign pk_rsp_dat_mergb[63:0] = _0197_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6062" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[31:30], 14'b00000000000000, img2sbuf_p0_rd_data[29:20], 6'b000000, img2sbuf_p0_rd_data[19:10], 6'b000000, img2sbuf_p0_rd_data[9:0], 6'b000000 };
  assign pk_rsp_dat_mergb[127:64] = _0199_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6064" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[63:62], 14'b00000000000000, img2sbuf_p0_rd_data[61:52], 6'b000000, img2sbuf_p0_rd_data[51:42], 6'b000000, img2sbuf_p0_rd_data[41:32], 6'b000000 };
  assign pk_rsp_dat_mergb[191:128] = _0201_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6066" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[95:94], 14'b00000000000000, img2sbuf_p0_rd_data[93:84], 6'b000000, img2sbuf_p0_rd_data[83:74], 6'b000000, img2sbuf_p0_rd_data[73:64], 6'b000000 };
  assign pk_rsp_dat_mergb[255:192] = _0203_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6068" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[127:126], 14'b00000000000000, img2sbuf_p0_rd_data[125:116], 6'b000000, img2sbuf_p0_rd_data[115:106], 6'b000000, img2sbuf_p0_rd_data[105:96], 6'b000000 };
  assign pk_rsp_dat_mergb[319:256] = _0205_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6070" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[159:158], 14'b00000000000000, img2sbuf_p0_rd_data[157:148], 6'b000000, img2sbuf_p0_rd_data[147:138], 6'b000000, img2sbuf_p0_rd_data[137:128], 6'b000000 };
  assign pk_rsp_dat_mergb[383:320] = _0207_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6072" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[191:190], 14'b00000000000000, img2sbuf_p0_rd_data[189:180], 6'b000000, img2sbuf_p0_rd_data[179:170], 6'b000000, img2sbuf_p0_rd_data[169:160], 6'b000000 };
  assign pk_rsp_dat_mergb[447:384] = _0209_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6074" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[223:222], 14'b00000000000000, img2sbuf_p0_rd_data[221:212], 6'b000000, img2sbuf_p0_rd_data[211:202], 6'b000000, img2sbuf_p0_rd_data[201:192], 6'b000000 };
  assign pk_rsp_dat_mergb[511:448] = _0211_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6076" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p0_rd_data[255:254], 14'b00000000000000, img2sbuf_p0_rd_data[253:244], 6'b000000, img2sbuf_p0_rd_data[243:234], 6'b000000, img2sbuf_p0_rd_data[233:224], 6'b000000 };
  assign pk_rsp_data_h1[63:0] = _0213_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6078" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[31:30], 14'b00000000000000, img2sbuf_p1_rd_data[29:20], 6'b000000, img2sbuf_p1_rd_data[19:10], 6'b000000, img2sbuf_p1_rd_data[9:0], 6'b000000 };
  assign pk_rsp_data_h1[127:64] = _0215_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6080" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[63:62], 14'b00000000000000, img2sbuf_p1_rd_data[61:52], 6'b000000, img2sbuf_p1_rd_data[51:42], 6'b000000, img2sbuf_p1_rd_data[41:32], 6'b000000 };
  assign pk_rsp_data_h1[191:128] = _0217_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6082" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[95:94], 14'b00000000000000, img2sbuf_p1_rd_data[93:84], 6'b000000, img2sbuf_p1_rd_data[83:74], 6'b000000, img2sbuf_p1_rd_data[73:64], 6'b000000 };
  assign pk_rsp_data_h1[255:192] = _0219_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6084" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[127:126], 14'b00000000000000, img2sbuf_p1_rd_data[125:116], 6'b000000, img2sbuf_p1_rd_data[115:106], 6'b000000, img2sbuf_p1_rd_data[105:96], 6'b000000 };
  assign pk_rsp_data_h1[319:256] = _0221_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6086" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[159:158], 14'b00000000000000, img2sbuf_p1_rd_data[157:148], 6'b000000, img2sbuf_p1_rd_data[147:138], 6'b000000, img2sbuf_p1_rd_data[137:128], 6'b000000 };
  assign pk_rsp_data_h1[383:320] = _0223_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6088" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[191:190], 14'b00000000000000, img2sbuf_p1_rd_data[189:180], 6'b000000, img2sbuf_p1_rd_data[179:170], 6'b000000, img2sbuf_p1_rd_data[169:160], 6'b000000 };
  assign pk_rsp_data_h1[447:384] = _0225_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6090" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[223:222], 14'b00000000000000, img2sbuf_p1_rd_data[221:212], 6'b000000, img2sbuf_p1_rd_data[211:202], 6'b000000, img2sbuf_p1_rd_data[201:192], 6'b000000 };
  assign pk_rsp_data_h1[511:448] = _0227_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6092" *) 64'b0000000000000000000000000000000000000000000000000000000000000000 : { img2sbuf_p1_rd_data[255:254], 14'b00000000000000, img2sbuf_p1_rd_data[253:244], 6'b000000, img2sbuf_p1_rd_data[243:234], 6'b000000, img2sbuf_p1_rd_data[233:224], 6'b000000 };
  assign pk_rsp_dat_mnorm[7:0] = _0229_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6101" *) 8'b00000000 : img2sbuf_p0_rd_data[7:0];
  assign pk_rsp_dat_mnorm[15:8] = _0231_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6103" *) 8'b00000000 : img2sbuf_p0_rd_data[15:8];
  assign pk_rsp_dat_mnorm[23:16] = _0233_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6105" *) 8'b00000000 : img2sbuf_p0_rd_data[23:16];
  assign pk_rsp_dat_mnorm[31:24] = _0235_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6107" *) 8'b00000000 : img2sbuf_p0_rd_data[31:24];
  assign pk_rsp_dat_mnorm[39:32] = _0237_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6109" *) 8'b00000000 : img2sbuf_p0_rd_data[39:32];
  assign pk_rsp_dat_mnorm[47:40] = _0239_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6111" *) 8'b00000000 : img2sbuf_p0_rd_data[47:40];
  assign pk_rsp_dat_mnorm[55:48] = _0241_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6113" *) 8'b00000000 : img2sbuf_p0_rd_data[55:48];
  assign pk_rsp_dat_mnorm[63:56] = _0243_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6115" *) 8'b00000000 : img2sbuf_p0_rd_data[63:56];
  assign pk_rsp_dat_mnorm[71:64] = _0245_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6117" *) 8'b00000000 : img2sbuf_p0_rd_data[71:64];
  assign pk_rsp_dat_mnorm[79:72] = _0247_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6119" *) 8'b00000000 : img2sbuf_p0_rd_data[79:72];
  assign pk_rsp_dat_mnorm[87:80] = _0249_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6121" *) 8'b00000000 : img2sbuf_p0_rd_data[87:80];
  assign pk_rsp_dat_mnorm[95:88] = _0251_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6123" *) 8'b00000000 : img2sbuf_p0_rd_data[95:88];
  assign pk_rsp_dat_mnorm[103:96] = _0253_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6125" *) 8'b00000000 : img2sbuf_p0_rd_data[103:96];
  assign pk_rsp_dat_mnorm[111:104] = _0255_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6127" *) 8'b00000000 : img2sbuf_p0_rd_data[111:104];
  assign pk_rsp_dat_mnorm[119:112] = _0257_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6129" *) 8'b00000000 : img2sbuf_p0_rd_data[119:112];
  assign pk_rsp_dat_mnorm[127:120] = _0259_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6131" *) 8'b00000000 : img2sbuf_p0_rd_data[127:120];
  assign pk_rsp_dat_mnorm[135:128] = _0261_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6133" *) 8'b00000000 : img2sbuf_p0_rd_data[135:128];
  assign pk_rsp_dat_mnorm[143:136] = _0263_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6135" *) 8'b00000000 : img2sbuf_p0_rd_data[143:136];
  assign pk_rsp_dat_mnorm[151:144] = _0265_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6137" *) 8'b00000000 : img2sbuf_p0_rd_data[151:144];
  assign pk_rsp_dat_mnorm[159:152] = _0267_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6139" *) 8'b00000000 : img2sbuf_p0_rd_data[159:152];
  assign pk_rsp_dat_mnorm[167:160] = _0269_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6141" *) 8'b00000000 : img2sbuf_p0_rd_data[167:160];
  assign pk_rsp_dat_mnorm[175:168] = _0271_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6143" *) 8'b00000000 : img2sbuf_p0_rd_data[175:168];
  assign pk_rsp_dat_mnorm[183:176] = _0273_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6145" *) 8'b00000000 : img2sbuf_p0_rd_data[183:176];
  assign pk_rsp_dat_mnorm[191:184] = _0275_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6147" *) 8'b00000000 : img2sbuf_p0_rd_data[191:184];
  assign pk_rsp_dat_mnorm[199:192] = _0277_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6149" *) 8'b00000000 : img2sbuf_p0_rd_data[199:192];
  assign pk_rsp_dat_mnorm[207:200] = _0279_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6151" *) 8'b00000000 : img2sbuf_p0_rd_data[207:200];
  assign pk_rsp_dat_mnorm[215:208] = _0281_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6153" *) 8'b00000000 : img2sbuf_p0_rd_data[215:208];
  assign pk_rsp_dat_mnorm[223:216] = _0283_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6155" *) 8'b00000000 : img2sbuf_p0_rd_data[223:216];
  assign pk_rsp_dat_mnorm[231:224] = _0285_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6157" *) 8'b00000000 : img2sbuf_p0_rd_data[231:224];
  assign pk_rsp_dat_mnorm[239:232] = _0287_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6159" *) 8'b00000000 : img2sbuf_p0_rd_data[239:232];
  assign pk_rsp_dat_mnorm[247:240] = _0289_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6161" *) 8'b00000000 : img2sbuf_p0_rd_data[247:240];
  assign pk_rsp_dat_mnorm[255:248] = _0291_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6163" *) 8'b00000000 : img2sbuf_p0_rd_data[255:248];
  assign pk_rsp_dat_mnorm[263:256] = _0293_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6165" *) 8'b00000000 : img2sbuf_p1_rd_data[7:0];
  assign pk_rsp_dat_mnorm[271:264] = _0295_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6167" *) 8'b00000000 : img2sbuf_p1_rd_data[15:8];
  assign pk_rsp_dat_mnorm[279:272] = _0297_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6169" *) 8'b00000000 : img2sbuf_p1_rd_data[23:16];
  assign pk_rsp_dat_mnorm[287:280] = _0299_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6171" *) 8'b00000000 : img2sbuf_p1_rd_data[31:24];
  assign pk_rsp_dat_mnorm[295:288] = _0301_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6173" *) 8'b00000000 : img2sbuf_p1_rd_data[39:32];
  assign pk_rsp_dat_mnorm[303:296] = _0303_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6175" *) 8'b00000000 : img2sbuf_p1_rd_data[47:40];
  assign pk_rsp_dat_mnorm[311:304] = _0305_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6177" *) 8'b00000000 : img2sbuf_p1_rd_data[55:48];
  assign pk_rsp_dat_mnorm[319:312] = _0307_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6179" *) 8'b00000000 : img2sbuf_p1_rd_data[63:56];
  assign pk_rsp_dat_mnorm[327:320] = _0309_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6181" *) 8'b00000000 : img2sbuf_p1_rd_data[71:64];
  assign pk_rsp_dat_mnorm[335:328] = _0311_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6183" *) 8'b00000000 : img2sbuf_p1_rd_data[79:72];
  assign pk_rsp_dat_mnorm[343:336] = _0313_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6185" *) 8'b00000000 : img2sbuf_p1_rd_data[87:80];
  assign pk_rsp_dat_mnorm[351:344] = _0315_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6187" *) 8'b00000000 : img2sbuf_p1_rd_data[95:88];
  assign pk_rsp_dat_mnorm[359:352] = _0317_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6189" *) 8'b00000000 : img2sbuf_p1_rd_data[103:96];
  assign pk_rsp_dat_mnorm[367:360] = _0319_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6191" *) 8'b00000000 : img2sbuf_p1_rd_data[111:104];
  assign pk_rsp_dat_mnorm[375:368] = _0321_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6193" *) 8'b00000000 : img2sbuf_p1_rd_data[119:112];
  assign pk_rsp_dat_mnorm[383:376] = _0323_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6195" *) 8'b00000000 : img2sbuf_p1_rd_data[127:120];
  assign pk_rsp_dat_mnorm[391:384] = _0325_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6197" *) 8'b00000000 : img2sbuf_p1_rd_data[135:128];
  assign pk_rsp_dat_mnorm[399:392] = _0327_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6199" *) 8'b00000000 : img2sbuf_p1_rd_data[143:136];
  assign pk_rsp_dat_mnorm[407:400] = _0329_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6201" *) 8'b00000000 : img2sbuf_p1_rd_data[151:144];
  assign pk_rsp_dat_mnorm[415:408] = _0331_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6203" *) 8'b00000000 : img2sbuf_p1_rd_data[159:152];
  assign pk_rsp_dat_mnorm[423:416] = _0333_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6205" *) 8'b00000000 : img2sbuf_p1_rd_data[167:160];
  assign pk_rsp_dat_mnorm[431:424] = _0335_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6207" *) 8'b00000000 : img2sbuf_p1_rd_data[175:168];
  assign pk_rsp_dat_mnorm[439:432] = _0337_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6209" *) 8'b00000000 : img2sbuf_p1_rd_data[183:176];
  assign pk_rsp_dat_mnorm[447:440] = _0339_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6211" *) 8'b00000000 : img2sbuf_p1_rd_data[191:184];
  assign pk_rsp_dat_mnorm[455:448] = _0341_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6213" *) 8'b00000000 : img2sbuf_p1_rd_data[199:192];
  assign pk_rsp_dat_mnorm[463:456] = _0343_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6215" *) 8'b00000000 : img2sbuf_p1_rd_data[207:200];
  assign pk_rsp_dat_mnorm[471:464] = _0345_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6217" *) 8'b00000000 : img2sbuf_p1_rd_data[215:208];
  assign pk_rsp_dat_mnorm[479:472] = _0347_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6219" *) 8'b00000000 : img2sbuf_p1_rd_data[223:216];
  assign pk_rsp_dat_mnorm[487:480] = _0349_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6221" *) 8'b00000000 : img2sbuf_p1_rd_data[231:224];
  assign pk_rsp_dat_mnorm[495:488] = _0351_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6223" *) 8'b00000000 : img2sbuf_p1_rd_data[239:232];
  assign pk_rsp_dat_mnorm[503:496] = _0353_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6225" *) 8'b00000000 : img2sbuf_p1_rd_data[247:240];
  assign pk_rsp_dat_mnorm[511:504] = _0355_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6227" *) 8'b00000000 : img2sbuf_p1_rd_data[255:248];
  assign dat_yuv[1519:0] = _0152_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6235" *) { pk_rsp_planar0_c0_d1[511:504], dat_l1_hi[495:480], pk_rsp_planar0_c0_d1[503:496], dat_l1_hi[479:464], pk_rsp_planar0_c0_d1[495:488], dat_l1_hi[463:448], pk_rsp_planar0_c0_d1[487:480], dat_l1_hi[447:432], pk_rsp_planar0_c0_d1[479:472], dat_l1_hi[431:416], pk_rsp_planar0_c0_d1[471:464], dat_l1_hi[415:400], pk_rsp_planar0_c0_d1[463:456], dat_l1_hi[399:384], pk_rsp_planar0_c0_d1[455:448], dat_l1_hi[383:368], pk_rsp_planar0_c0_d1[447:440], dat_l1_hi[367:352], pk_rsp_planar0_c0_d1[439:432], dat_l1_hi[351:336], pk_rsp_planar0_c0_d1[431:424], dat_l1_hi[335:320], pk_rsp_planar0_c0_d1[423:416], dat_l1_hi[319:304], pk_rsp_planar0_c0_d1[415:408], dat_l1_hi[303:288], pk_rsp_planar0_c0_d1[407:400], dat_l1_hi[287:272], pk_rsp_planar0_c0_d1[399:392], dat_l1_hi[271:256], pk_rsp_planar0_c0_d1[391:384], dat_l1_hi[255:240], pk_rsp_planar0_c0_d1[383:376], dat_l1_hi[239:224], pk_rsp_planar0_c0_d1[375:368], dat_l1_hi[223:208], pk_rsp_planar0_c0_d1[367:360], dat_l1_hi[207:192], pk_rsp_planar0_c0_d1[359:352], dat_l1_hi[191:176], pk_rsp_planar0_c0_d1[351:344], dat_l1_hi[175:160], pk_rsp_planar0_c0_d1[343:336], dat_l1_hi[159:144], pk_rsp_planar0_c0_d1[335:328], dat_l1_hi[143:128], pk_rsp_planar0_c0_d1[327:320], dat_l1_hi[127:112], pk_rsp_planar0_c0_d1[319:312], dat_l1_hi[111:96], pk_rsp_planar0_c0_d1[311:304], dat_l1_hi[95:80], pk_rsp_planar0_c0_d1[303:296], dat_l1_hi[79:64], pk_rsp_planar0_c0_d1[295:288], dat_l1_hi[63:48], pk_rsp_planar0_c0_d1[287:280], dat_l1_hi[47:32], pk_rsp_planar0_c0_d1[279:272], dat_l1_hi[31:16], pk_rsp_planar0_c0_d1[271:264], dat_l1_hi[15:0], pk_rsp_planar0_c0_d1[263:256], dat_l1_lo[511:496], pk_rsp_planar0_c0_d1[255:248], dat_l1_lo[495:480], pk_rsp_planar0_c0_d1[247:240], dat_l1_lo[479:464], pk_rsp_planar0_c0_d1[239:232], dat_l1_lo[463:448], pk_rsp_planar0_c0_d1[231:224], dat_l1_lo[447:432], pk_rsp_planar0_c0_d1[223:216], dat_l1_lo[431:416], pk_rsp_planar0_c0_d1[215:208], dat_l1_lo[415:400], pk_rsp_planar0_c0_d1[207:200], dat_l1_lo[399:384], pk_rsp_planar0_c0_d1[199:192], dat_l1_lo[383:368], pk_rsp_planar0_c0_d1[191:184], dat_l1_lo[367:352], pk_rsp_planar0_c0_d1[183:176], dat_l1_lo[351:336], pk_rsp_planar0_c0_d1[175:168], dat_l1_lo[335:320], pk_rsp_planar0_c0_d1[167:160], dat_l1_lo[319:304], pk_rsp_planar0_c0_d1[159:152], dat_l1_lo[303:288], pk_rsp_planar0_c0_d1[151:144], dat_l1_lo[287:272], pk_rsp_planar0_c0_d1[143:136], dat_l1_lo[271:256], pk_rsp_planar0_c0_d1[135:128], dat_l1_lo[255:240], pk_rsp_planar0_c0_d1[127:120], dat_l1_lo[239:224], pk_rsp_planar0_c0_d1[119:112], dat_l1_lo[223:208], pk_rsp_planar0_c0_d1[111:104], dat_l1_lo[207:192], pk_rsp_planar0_c0_d1[103:96], dat_l1_lo[191:176], pk_rsp_planar0_c0_d1[95:88], dat_l1_lo[175:160], pk_rsp_planar0_c0_d1[87:80], dat_l1_lo[159:144], pk_rsp_planar0_c0_d1[79:72], dat_l1_lo[143:128], pk_rsp_planar0_c0_d1[71:64], dat_l1_lo[127:112], pk_rsp_planar0_c0_d1[63:56], dat_l1_lo[111:96], pk_rsp_planar0_c0_d1[55:48], dat_l1_lo[95:80], pk_rsp_planar0_c0_d1[47:40], dat_l1_lo[79:64], pk_rsp_planar0_c0_d1[39:32], dat_l1_lo[63:48], pk_rsp_planar0_c0_d1[31:24], dat_l1_lo[47:32], pk_rsp_planar0_c0_d1[23:16], dat_l1_lo[31:16], pk_rsp_planar0_c0_d1[15:8], dat_l1_lo[15:0], pk_rsp_planar0_c0_d1[7:0] } : { dat_l1_hi[495:480], pk_rsp_planar0_c0_d1[511:496], dat_l1_hi[479:448], pk_rsp_planar0_c0_d1[495:480], dat_l1_hi[447:416], pk_rsp_planar0_c0_d1[479:464], dat_l1_hi[415:384], pk_rsp_planar0_c0_d1[463:448], dat_l1_hi[383:352], pk_rsp_planar0_c0_d1[447:432], dat_l1_hi[351:320], pk_rsp_planar0_c0_d1[431:416], dat_l1_hi[319:288], pk_rsp_planar0_c0_d1[415:400], dat_l1_hi[287:256], pk_rsp_planar0_c0_d1[399:384], dat_l1_hi[255:224], pk_rsp_planar0_c0_d1[383:368], dat_l1_hi[223:192], pk_rsp_planar0_c0_d1[367:352], dat_l1_hi[191:160], pk_rsp_planar0_c0_d1[351:336], dat_l1_hi[159:128], pk_rsp_planar0_c0_d1[335:320], dat_l1_hi[127:96], pk_rsp_planar0_c0_d1[319:304], dat_l1_hi[95:64], pk_rsp_planar0_c0_d1[303:288], dat_l1_hi[63:32], pk_rsp_planar0_c0_d1[287:272], dat_l1_hi[31:0], pk_rsp_planar0_c0_d1[271:256], dat_l1_lo[511:480], pk_rsp_planar0_c0_d1[255:240], dat_l1_lo[479:448], pk_rsp_planar0_c0_d1[239:224], dat_l1_lo[447:416], pk_rsp_planar0_c0_d1[223:208], dat_l1_lo[415:384], pk_rsp_planar0_c0_d1[207:192], dat_l1_lo[383:352], pk_rsp_planar0_c0_d1[191:176], dat_l1_lo[351:320], pk_rsp_planar0_c0_d1[175:160], dat_l1_lo[319:288], pk_rsp_planar0_c0_d1[159:144], dat_l1_lo[287:256], pk_rsp_planar0_c0_d1[143:128], dat_l1_lo[255:224], pk_rsp_planar0_c0_d1[127:112], dat_l1_lo[223:192], pk_rsp_planar0_c0_d1[111:96], dat_l1_lo[191:160], pk_rsp_planar0_c0_d1[95:80], dat_l1_lo[159:128], pk_rsp_planar0_c0_d1[79:64], dat_l1_lo[127:96], pk_rsp_planar0_c0_d1[63:48], dat_l1_lo[95:64], pk_rsp_planar0_c0_d1[47:32], dat_l1_lo[63:32], pk_rsp_planar0_c0_d1[31:16], dat_l1_lo[31:0], pk_rsp_planar0_c0_d1[15:0] };
  assign pad_mask_yuv[189:0] = _0152_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6272" *) { mask_pad_planar0_c0_d1[63], pad_mask_l1_hi[61:60], mask_pad_planar0_c0_d1[62], pad_mask_l1_hi[59:58], mask_pad_planar0_c0_d1[61], pad_mask_l1_hi[57:56], mask_pad_planar0_c0_d1[60], pad_mask_l1_hi[55:54], mask_pad_planar0_c0_d1[59], pad_mask_l1_hi[53:52], mask_pad_planar0_c0_d1[58], pad_mask_l1_hi[51:50], mask_pad_planar0_c0_d1[57], pad_mask_l1_hi[49:48], mask_pad_planar0_c0_d1[56], pad_mask_l1_hi[47:46], mask_pad_planar0_c0_d1[55], pad_mask_l1_hi[45:44], mask_pad_planar0_c0_d1[54], pad_mask_l1_hi[43:42], mask_pad_planar0_c0_d1[53], pad_mask_l1_hi[41:40], mask_pad_planar0_c0_d1[52], pad_mask_l1_hi[39:38], mask_pad_planar0_c0_d1[51], pad_mask_l1_hi[37:36], mask_pad_planar0_c0_d1[50], pad_mask_l1_hi[35:34], mask_pad_planar0_c0_d1[49], pad_mask_l1_hi[33:32], mask_pad_planar0_c0_d1[48], pad_mask_l1_hi[31:30], mask_pad_planar0_c0_d1[47], pad_mask_l1_hi[29:28], mask_pad_planar0_c0_d1[46], pad_mask_l1_hi[27:26], mask_pad_planar0_c0_d1[45], pad_mask_l1_hi[25:24], mask_pad_planar0_c0_d1[44], pad_mask_l1_hi[23:22], mask_pad_planar0_c0_d1[43], pad_mask_l1_hi[21:20], mask_pad_planar0_c0_d1[42], pad_mask_l1_hi[19:18], mask_pad_planar0_c0_d1[41], pad_mask_l1_hi[17:16], mask_pad_planar0_c0_d1[40], pad_mask_l1_hi[15:14], mask_pad_planar0_c0_d1[39], pad_mask_l1_hi[13:12], mask_pad_planar0_c0_d1[38], pad_mask_l1_hi[11:10], mask_pad_planar0_c0_d1[37], pad_mask_l1_hi[9:8], mask_pad_planar0_c0_d1[36], pad_mask_l1_hi[7:6], mask_pad_planar0_c0_d1[35], pad_mask_l1_hi[5:4], mask_pad_planar0_c0_d1[34], pad_mask_l1_hi[3:2], mask_pad_planar0_c0_d1[33], pad_mask_l1_hi[1:0], mask_pad_planar0_c0_d1[32], pad_mask_l1_lo[63:62], mask_pad_planar0_c0_d1[31], pad_mask_l1_lo[61:60], mask_pad_planar0_c0_d1[30], pad_mask_l1_lo[59:58], mask_pad_planar0_c0_d1[29], pad_mask_l1_lo[57:56], mask_pad_planar0_c0_d1[28], pad_mask_l1_lo[55:54], mask_pad_planar0_c0_d1[27], pad_mask_l1_lo[53:52], mask_pad_planar0_c0_d1[26], pad_mask_l1_lo[51:50], mask_pad_planar0_c0_d1[25], pad_mask_l1_lo[49:48], mask_pad_planar0_c0_d1[24], pad_mask_l1_lo[47:46], mask_pad_planar0_c0_d1[23], pad_mask_l1_lo[45:44], mask_pad_planar0_c0_d1[22], pad_mask_l1_lo[43:42], mask_pad_planar0_c0_d1[21], pad_mask_l1_lo[41:40], mask_pad_planar0_c0_d1[20], pad_mask_l1_lo[39:38], mask_pad_planar0_c0_d1[19], pad_mask_l1_lo[37:36], mask_pad_planar0_c0_d1[18], pad_mask_l1_lo[35:34], mask_pad_planar0_c0_d1[17], pad_mask_l1_lo[33:32], mask_pad_planar0_c0_d1[16], pad_mask_l1_lo[31:30], mask_pad_planar0_c0_d1[15], pad_mask_l1_lo[29:28], mask_pad_planar0_c0_d1[14], pad_mask_l1_lo[27:26], mask_pad_planar0_c0_d1[13], pad_mask_l1_lo[25:24], mask_pad_planar0_c0_d1[12], pad_mask_l1_lo[23:22], mask_pad_planar0_c0_d1[11], pad_mask_l1_lo[21:20], mask_pad_planar0_c0_d1[10], pad_mask_l1_lo[19:18], mask_pad_planar0_c0_d1[9], pad_mask_l1_lo[17:16], mask_pad_planar0_c0_d1[8], pad_mask_l1_lo[15:14], mask_pad_planar0_c0_d1[7], pad_mask_l1_lo[13:12], mask_pad_planar0_c0_d1[6], pad_mask_l1_lo[11:10], mask_pad_planar0_c0_d1[5], pad_mask_l1_lo[9:8], mask_pad_planar0_c0_d1[4], pad_mask_l1_lo[7:6], mask_pad_planar0_c0_d1[3], pad_mask_l1_lo[5:4], mask_pad_planar0_c0_d1[2], pad_mask_l1_lo[3:2], mask_pad_planar0_c0_d1[1], pad_mask_l1_lo[1:0], mask_pad_planar0_c0_d1[0] } : { pad_mask_l1_hi[61:60], mask_pad_planar0_c0_d1[63:62], pad_mask_l1_hi[59:56], mask_pad_planar0_c0_d1[61:60], pad_mask_l1_hi[55:52], mask_pad_planar0_c0_d1[59:58], pad_mask_l1_hi[51:48], mask_pad_planar0_c0_d1[57:56], pad_mask_l1_hi[47:44], mask_pad_planar0_c0_d1[55:54], pad_mask_l1_hi[43:40], mask_pad_planar0_c0_d1[53:52], pad_mask_l1_hi[39:36], mask_pad_planar0_c0_d1[51:50], pad_mask_l1_hi[35:32], mask_pad_planar0_c0_d1[49:48], pad_mask_l1_hi[31:28], mask_pad_planar0_c0_d1[47:46], pad_mask_l1_hi[27:24], mask_pad_planar0_c0_d1[45:44], pad_mask_l1_hi[23:20], mask_pad_planar0_c0_d1[43:42], pad_mask_l1_hi[19:16], mask_pad_planar0_c0_d1[41:40], pad_mask_l1_hi[15:12], mask_pad_planar0_c0_d1[39:38], pad_mask_l1_hi[11:8], mask_pad_planar0_c0_d1[37:36], pad_mask_l1_hi[7:4], mask_pad_planar0_c0_d1[35:34], pad_mask_l1_hi[3:0], mask_pad_planar0_c0_d1[33:32], pad_mask_l1_lo[63:60], mask_pad_planar0_c0_d1[31:30], pad_mask_l1_lo[59:56], mask_pad_planar0_c0_d1[29:28], pad_mask_l1_lo[55:52], mask_pad_planar0_c0_d1[27:26], pad_mask_l1_lo[51:48], mask_pad_planar0_c0_d1[25:24], pad_mask_l1_lo[47:44], mask_pad_planar0_c0_d1[23:22], pad_mask_l1_lo[43:40], mask_pad_planar0_c0_d1[21:20], pad_mask_l1_lo[39:36], mask_pad_planar0_c0_d1[19:18], pad_mask_l1_lo[35:32], mask_pad_planar0_c0_d1[17:16], pad_mask_l1_lo[31:28], mask_pad_planar0_c0_d1[15:14], pad_mask_l1_lo[27:24], mask_pad_planar0_c0_d1[13:12], pad_mask_l1_lo[23:20], mask_pad_planar0_c0_d1[11:10], pad_mask_l1_lo[19:16], mask_pad_planar0_c0_d1[9:8], pad_mask_l1_lo[15:12], mask_pad_planar0_c0_d1[7:6], pad_mask_l1_lo[11:8], mask_pad_planar0_c0_d1[5:4], pad_mask_l1_lo[7:4], mask_pad_planar0_c0_d1[3:2], pad_mask_l1_lo[3:0], mask_pad_planar0_c0_d1[1:0] };
  assign pk_rsp_pad_mask_h1 = pixel_packed_10b ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6277" *) { rd_p1_pad_mask_d3[31], rd_p1_pad_mask_d3[31:30], rd_p1_pad_mask_d3[30:29], rd_p1_pad_mask_d3[29:28], rd_p1_pad_mask_d3[28:27], rd_p1_pad_mask_d3[27:26], rd_p1_pad_mask_d3[26:25], rd_p1_pad_mask_d3[25:24], rd_p1_pad_mask_d3[24:23], rd_p1_pad_mask_d3[23:22], rd_p1_pad_mask_d3[22:21], rd_p1_pad_mask_d3[21:20], rd_p1_pad_mask_d3[20:19], rd_p1_pad_mask_d3[19:18], rd_p1_pad_mask_d3[18:17], rd_p1_pad_mask_d3[17:16], rd_p1_pad_mask_d3[16:15], rd_p1_pad_mask_d3[15:14], rd_p1_pad_mask_d3[14:13], rd_p1_pad_mask_d3[13:12], rd_p1_pad_mask_d3[12:11], rd_p1_pad_mask_d3[11:10], rd_p1_pad_mask_d3[10:9], rd_p1_pad_mask_d3[9:8], rd_p1_pad_mask_d3[8:7], rd_p1_pad_mask_d3[7:6], rd_p1_pad_mask_d3[6:5], rd_p1_pad_mask_d3[5:4], rd_p1_pad_mask_d3[4:3], rd_p1_pad_mask_d3[3:2], rd_p1_pad_mask_d3[2:1], rd_p1_pad_mask_d3[1:0], rd_p1_pad_mask_d3[0] } : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign mn_ch1_4 = _0374_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6817" *) { reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry } : { reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry };
  assign mn_16b_mnorm[15:0] = rd_p0_zero_mask_d3[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6822" *) 16'b0000000000000000 : mn_ch1_4[15:0];
  assign mn_8b_mnorm[31:16] = rd_p0_zero_mask_d3[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6823" *) 16'b0000000000000000 : mn_ch1_4[31:16];
  assign mn_8b_mnorm[47:32] = rd_p0_zero_mask_d3[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6824" *) 16'b0000000000000000 : mn_ch1_4[47:32];
  assign mn_8b_mnorm[63:48] = rd_p0_zero_mask_d3[3] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6825" *) 16'b0000000000000000 : mn_ch1_4[63:48];
  assign mn_8b_mnorm[79:64] = rd_p0_zero_mask_d3[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6826" *) 16'b0000000000000000 : mn_ch1_4[79:64];
  assign mn_8b_mnorm[95:80] = rd_p0_zero_mask_d3[5] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6827" *) 16'b0000000000000000 : mn_ch1_4[95:80];
  assign mn_8b_mnorm[111:96] = rd_p0_zero_mask_d3[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6828" *) 16'b0000000000000000 : mn_ch1_4[111:96];
  assign mn_8b_mnorm[127:112] = rd_p0_zero_mask_d3[7] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6829" *) 16'b0000000000000000 : mn_ch1_4[127:112];
  assign mn_8b_mnorm[143:128] = rd_p0_zero_mask_d3[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6830" *) 16'b0000000000000000 : mn_ch1_4[143:128];
  assign mn_8b_mnorm[159:144] = rd_p0_zero_mask_d3[9] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6831" *) 16'b0000000000000000 : mn_ch1_4[159:144];
  assign mn_8b_mnorm[175:160] = rd_p0_zero_mask_d3[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6832" *) 16'b0000000000000000 : mn_ch1_4[175:160];
  assign mn_8b_mnorm[191:176] = rd_p0_zero_mask_d3[11] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6833" *) 16'b0000000000000000 : mn_ch1_4[191:176];
  assign mn_8b_mnorm[207:192] = rd_p0_zero_mask_d3[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6834" *) 16'b0000000000000000 : mn_ch1_4[207:192];
  assign mn_8b_mnorm[223:208] = rd_p0_zero_mask_d3[13] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6835" *) 16'b0000000000000000 : mn_ch1_4[223:208];
  assign mn_8b_mnorm[239:224] = rd_p0_zero_mask_d3[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6836" *) 16'b0000000000000000 : mn_ch1_4[239:224];
  assign mn_8b_mnorm[255:240] = rd_p0_zero_mask_d3[15] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6837" *) 16'b0000000000000000 : mn_ch1_4[255:240];
  assign mn_8b_mnorm[271:256] = rd_p0_zero_mask_d3[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6838" *) 16'b0000000000000000 : mn_ch1_4[271:256];
  assign mn_8b_mnorm[287:272] = rd_p0_zero_mask_d3[17] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6839" *) 16'b0000000000000000 : mn_ch1_4[287:272];
  assign mn_8b_mnorm[303:288] = rd_p0_zero_mask_d3[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6840" *) 16'b0000000000000000 : mn_ch1_4[303:288];
  assign mn_8b_mnorm[319:304] = rd_p0_zero_mask_d3[19] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6841" *) 16'b0000000000000000 : mn_ch1_4[319:304];
  assign mn_8b_mnorm[335:320] = rd_p0_zero_mask_d3[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6842" *) 16'b0000000000000000 : mn_ch1_4[335:320];
  assign mn_8b_mnorm[351:336] = rd_p0_zero_mask_d3[21] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6843" *) 16'b0000000000000000 : mn_ch1_4[351:336];
  assign mn_8b_mnorm[367:352] = rd_p0_zero_mask_d3[22] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6844" *) 16'b0000000000000000 : mn_ch1_4[367:352];
  assign mn_8b_mnorm[383:368] = rd_p0_zero_mask_d3[23] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6845" *) 16'b0000000000000000 : mn_ch1_4[383:368];
  assign mn_8b_mnorm[399:384] = rd_p0_zero_mask_d3[24] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6846" *) 16'b0000000000000000 : mn_ch1_4[399:384];
  assign mn_8b_mnorm[415:400] = rd_p0_zero_mask_d3[25] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6847" *) 16'b0000000000000000 : mn_ch1_4[415:400];
  assign mn_8b_mnorm[431:416] = rd_p0_zero_mask_d3[26] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6848" *) 16'b0000000000000000 : mn_ch1_4[431:416];
  assign mn_8b_mnorm[447:432] = rd_p0_zero_mask_d3[27] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6849" *) 16'b0000000000000000 : mn_ch1_4[447:432];
  assign mn_8b_mnorm[463:448] = rd_p0_zero_mask_d3[28] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6850" *) 16'b0000000000000000 : mn_ch1_4[463:448];
  assign mn_8b_mnorm[479:464] = rd_p0_zero_mask_d3[29] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6851" *) 16'b0000000000000000 : mn_ch1_4[479:464];
  assign mn_8b_mnorm[495:480] = rd_p0_zero_mask_d3[30] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6852" *) 16'b0000000000000000 : mn_ch1_4[495:480];
  assign mn_8b_mnorm[511:496] = rd_p0_zero_mask_d3[31] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6853" *) 16'b0000000000000000 : mn_ch1_4[511:496];
  assign mn_8b_mnorm[527:512] = rd_p1_zero_mask_d3[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6854" *) 16'b0000000000000000 : mn_ch1_4[527:512];
  assign mn_8b_mnorm[543:528] = rd_p1_zero_mask_d3[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6855" *) 16'b0000000000000000 : mn_ch1_4[543:528];
  assign mn_8b_mnorm[559:544] = rd_p1_zero_mask_d3[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6856" *) 16'b0000000000000000 : mn_ch1_4[559:544];
  assign mn_8b_mnorm[575:560] = rd_p1_zero_mask_d3[3] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6857" *) 16'b0000000000000000 : mn_ch1_4[575:560];
  assign mn_8b_mnorm[591:576] = rd_p1_zero_mask_d3[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6858" *) 16'b0000000000000000 : mn_ch1_4[591:576];
  assign mn_8b_mnorm[607:592] = rd_p1_zero_mask_d3[5] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6859" *) 16'b0000000000000000 : mn_ch1_4[607:592];
  assign mn_8b_mnorm[623:608] = rd_p1_zero_mask_d3[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6860" *) 16'b0000000000000000 : mn_ch1_4[623:608];
  assign mn_8b_mnorm[639:624] = rd_p1_zero_mask_d3[7] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6861" *) 16'b0000000000000000 : mn_ch1_4[639:624];
  assign mn_8b_mnorm[655:640] = rd_p1_zero_mask_d3[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6862" *) 16'b0000000000000000 : mn_ch1_4[655:640];
  assign mn_8b_mnorm[671:656] = rd_p1_zero_mask_d3[9] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6863" *) 16'b0000000000000000 : mn_ch1_4[671:656];
  assign mn_8b_mnorm[687:672] = rd_p1_zero_mask_d3[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6864" *) 16'b0000000000000000 : mn_ch1_4[687:672];
  assign mn_8b_mnorm[703:688] = rd_p1_zero_mask_d3[11] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6865" *) 16'b0000000000000000 : mn_ch1_4[703:688];
  assign mn_8b_mnorm[719:704] = rd_p1_zero_mask_d3[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6866" *) 16'b0000000000000000 : mn_ch1_4[719:704];
  assign mn_8b_mnorm[735:720] = rd_p1_zero_mask_d3[13] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6867" *) 16'b0000000000000000 : mn_ch1_4[735:720];
  assign mn_8b_mnorm[751:736] = rd_p1_zero_mask_d3[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6868" *) 16'b0000000000000000 : mn_ch1_4[751:736];
  assign mn_8b_mnorm[767:752] = rd_p1_zero_mask_d3[15] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6869" *) 16'b0000000000000000 : mn_ch1_4[767:752];
  assign mn_8b_mnorm[783:768] = rd_p1_zero_mask_d3[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6870" *) 16'b0000000000000000 : mn_ch1_4[783:768];
  assign mn_8b_mnorm[799:784] = rd_p1_zero_mask_d3[17] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6871" *) 16'b0000000000000000 : mn_ch1_4[799:784];
  assign mn_8b_mnorm[815:800] = rd_p1_zero_mask_d3[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6872" *) 16'b0000000000000000 : mn_ch1_4[815:800];
  assign mn_8b_mnorm[831:816] = rd_p1_zero_mask_d3[19] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6873" *) 16'b0000000000000000 : mn_ch1_4[831:816];
  assign mn_8b_mnorm[847:832] = rd_p1_zero_mask_d3[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6874" *) 16'b0000000000000000 : mn_ch1_4[847:832];
  assign mn_8b_mnorm[863:848] = rd_p1_zero_mask_d3[21] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6875" *) 16'b0000000000000000 : mn_ch1_4[863:848];
  assign mn_8b_mnorm[879:864] = rd_p1_zero_mask_d3[22] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6876" *) 16'b0000000000000000 : mn_ch1_4[879:864];
  assign mn_8b_mnorm[895:880] = rd_p1_zero_mask_d3[23] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6877" *) 16'b0000000000000000 : mn_ch1_4[895:880];
  assign mn_8b_mnorm[911:896] = rd_p1_zero_mask_d3[24] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6878" *) 16'b0000000000000000 : mn_ch1_4[911:896];
  assign mn_8b_mnorm[927:912] = rd_p1_zero_mask_d3[25] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6879" *) 16'b0000000000000000 : mn_ch1_4[927:912];
  assign mn_8b_mnorm[943:928] = rd_p1_zero_mask_d3[26] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6880" *) 16'b0000000000000000 : mn_ch1_4[943:928];
  assign mn_8b_mnorm[959:944] = rd_p1_zero_mask_d3[27] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6881" *) 16'b0000000000000000 : mn_ch1_4[959:944];
  assign mn_8b_mnorm[975:960] = rd_p1_zero_mask_d3[28] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6882" *) 16'b0000000000000000 : mn_ch1_4[975:960];
  assign mn_8b_mnorm[991:976] = rd_p1_zero_mask_d3[29] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6883" *) 16'b0000000000000000 : mn_ch1_4[991:976];
  assign mn_8b_mnorm[1007:992] = rd_p1_zero_mask_d3[30] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6884" *) 16'b0000000000000000 : mn_ch1_4[1007:992];
  assign mn_8b_mnorm[1023:1008] = rd_p1_zero_mask_d3[31] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6885" *) 16'b0000000000000000 : mn_ch1_4[1023:1008];
  assign mn_16b_mnorm[31:16] = rd_p0_zero_mask_d3[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6892" *) 16'b0000000000000000 : mn_ch1_4[31:16];
  assign mn_16b_mnorm[47:32] = rd_p0_zero_mask_d3[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6893" *) 16'b0000000000000000 : mn_ch1_4[47:32];
  assign mn_16b_mnorm[63:48] = rd_p0_zero_mask_d3[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6894" *) 16'b0000000000000000 : mn_ch1_4[63:48];
  assign mn_16b_mnorm[79:64] = rd_p0_zero_mask_d3[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6895" *) 16'b0000000000000000 : mn_ch1_4[79:64];
  assign mn_16b_mnorm[95:80] = rd_p0_zero_mask_d3[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6896" *) 16'b0000000000000000 : mn_ch1_4[95:80];
  assign mn_16b_mnorm[111:96] = rd_p0_zero_mask_d3[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6897" *) 16'b0000000000000000 : mn_ch1_4[111:96];
  assign mn_16b_mnorm[127:112] = rd_p0_zero_mask_d3[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6898" *) 16'b0000000000000000 : mn_ch1_4[127:112];
  assign mn_16b_mnorm[143:128] = rd_p0_zero_mask_d3[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6899" *) 16'b0000000000000000 : mn_ch1_4[143:128];
  assign mn_16b_mnorm[159:144] = rd_p0_zero_mask_d3[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6900" *) 16'b0000000000000000 : mn_ch1_4[159:144];
  assign mn_16b_mnorm[175:160] = rd_p0_zero_mask_d3[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6901" *) 16'b0000000000000000 : mn_ch1_4[175:160];
  assign mn_16b_mnorm[191:176] = rd_p0_zero_mask_d3[22] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6902" *) 16'b0000000000000000 : mn_ch1_4[191:176];
  assign mn_16b_mnorm[207:192] = rd_p0_zero_mask_d3[24] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6903" *) 16'b0000000000000000 : mn_ch1_4[207:192];
  assign mn_16b_mnorm[223:208] = rd_p0_zero_mask_d3[26] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6904" *) 16'b0000000000000000 : mn_ch1_4[223:208];
  assign mn_16b_mnorm[239:224] = rd_p0_zero_mask_d3[28] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6905" *) 16'b0000000000000000 : mn_ch1_4[239:224];
  assign mn_16b_mnorm[255:240] = rd_p0_zero_mask_d3[30] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6906" *) 16'b0000000000000000 : mn_ch1_4[255:240];
  assign mn_16b_mnorm[271:256] = rd_p1_zero_mask_d3[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6907" *) 16'b0000000000000000 : mn_ch1_4[271:256];
  assign mn_16b_mnorm[287:272] = rd_p1_zero_mask_d3[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6908" *) 16'b0000000000000000 : mn_ch1_4[287:272];
  assign mn_16b_mnorm[303:288] = rd_p1_zero_mask_d3[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6909" *) 16'b0000000000000000 : mn_ch1_4[303:288];
  assign mn_16b_mnorm[319:304] = rd_p1_zero_mask_d3[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6910" *) 16'b0000000000000000 : mn_ch1_4[319:304];
  assign mn_16b_mnorm[335:320] = rd_p1_zero_mask_d3[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6911" *) 16'b0000000000000000 : mn_ch1_4[335:320];
  assign mn_16b_mnorm[351:336] = rd_p1_zero_mask_d3[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6912" *) 16'b0000000000000000 : mn_ch1_4[351:336];
  assign mn_16b_mnorm[367:352] = rd_p1_zero_mask_d3[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6913" *) 16'b0000000000000000 : mn_ch1_4[367:352];
  assign mn_16b_mnorm[383:368] = rd_p1_zero_mask_d3[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6914" *) 16'b0000000000000000 : mn_ch1_4[383:368];
  assign mn_16b_mnorm[399:384] = rd_p1_zero_mask_d3[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6915" *) 16'b0000000000000000 : mn_ch1_4[399:384];
  assign mn_16b_mnorm[415:400] = rd_p1_zero_mask_d3[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6916" *) 16'b0000000000000000 : mn_ch1_4[415:400];
  assign mn_16b_mnorm[431:416] = rd_p1_zero_mask_d3[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6917" *) 16'b0000000000000000 : mn_ch1_4[431:416];
  assign mn_16b_mnorm[447:432] = rd_p1_zero_mask_d3[22] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6918" *) 16'b0000000000000000 : mn_ch1_4[447:432];
  assign mn_16b_mnorm[463:448] = rd_p1_zero_mask_d3[24] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6919" *) 16'b0000000000000000 : mn_ch1_4[463:448];
  assign mn_16b_mnorm[479:464] = rd_p1_zero_mask_d3[26] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6920" *) 16'b0000000000000000 : mn_ch1_4[479:464];
  assign mn_16b_mnorm[495:480] = rd_p1_zero_mask_d3[28] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6921" *) 16'b0000000000000000 : mn_ch1_4[495:480];
  assign mn_16b_mnorm[511:496] = rd_p1_zero_mask_d3[30] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6922" *) 16'b0000000000000000 : mn_ch1_4[511:496];
  assign mn_16b_myuv[47:0] = mn_mask_y_d1[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6928" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[95:48] = mn_mask_y_d1[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6929" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[95:48] = mn_mask_uv_lo[0] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6930" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[191:144] = mn_mask_uv_lo[1] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6931" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[143:96] = mn_mask_uv_lo[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6932" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[287:240] = mn_mask_uv_lo[3] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6933" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[191:144] = mn_mask_y_d1[2] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6934" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[383:336] = mn_mask_y_d1[3] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6935" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[239:192] = mn_mask_uv_lo[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6936" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[479:432] = mn_mask_uv_lo[5] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6937" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[287:240] = mn_mask_uv_lo[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6938" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[575:528] = mn_mask_uv_lo[7] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6939" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[335:288] = mn_mask_y_d1[4] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6940" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[671:624] = mn_mask_y_d1[5] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6941" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[383:336] = mn_mask_uv_lo[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6942" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[767:720] = mn_mask_uv_lo[9] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6943" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[431:384] = mn_mask_uv_lo[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6944" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[863:816] = mn_mask_uv_lo[11] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6945" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[479:432] = mn_mask_y_d1[6] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6946" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[959:912] = mn_mask_y_d1[7] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6947" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[527:480] = mn_mask_uv_lo[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6948" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1055:1008] = mn_mask_uv_lo[13] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6949" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[575:528] = mn_mask_uv_lo[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6950" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1151:1104] = mn_mask_uv_lo[15] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6951" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[623:576] = mn_mask_y_d1[8] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6952" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1247:1200] = mn_mask_y_d1[9] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6953" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[671:624] = mn_mask_uv_lo[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6954" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1343:1296] = mn_mask_uv_lo[17] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6955" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[719:672] = mn_mask_uv_lo[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6956" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1439:1392] = mn_mask_uv_lo[19] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6957" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[767:720] = mn_mask_y_d1[10] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6958" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1535:1488] = mn_mask_y_d1[11] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6959" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[815:768] = mn_mask_uv_lo[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6960" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1631:1584] = mn_mask_uv_lo[21] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6961" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[863:816] = mn_mask_uv_lo[22] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6962" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1727:1680] = mn_mask_uv_lo[23] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6963" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[911:864] = mn_mask_y_d1[12] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6964" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1823:1776] = mn_mask_y_d1[13] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6965" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[959:912] = mn_mask_uv_lo[24] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6966" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[1919:1872] = mn_mask_uv_lo[25] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6967" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1007:960] = mn_mask_uv_lo[26] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6968" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2015:1968] = mn_mask_uv_lo[27] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6969" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1055:1008] = mn_mask_y_d1[14] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6970" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2111:2064] = mn_mask_y_d1[15] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6971" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1103:1056] = mn_mask_uv_lo[28] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6972" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2207:2160] = mn_mask_uv_lo[29] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6973" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1151:1104] = mn_mask_uv_lo[30] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6974" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2303:2256] = mn_mask_uv_lo[31] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6975" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1199:1152] = mn_mask_y_d1[16] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6976" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2399:2352] = mn_mask_y_d1[17] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6977" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1247:1200] = mn_mask_uv_lo[32] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6978" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2495:2448] = mn_mask_uv_lo[33] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6979" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1295:1248] = mn_mask_uv_lo[34] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6980" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2591:2544] = mn_mask_uv_lo[35] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6981" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1343:1296] = mn_mask_y_d1[18] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6982" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2687:2640] = mn_mask_y_d1[19] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6983" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1391:1344] = mn_mask_uv_lo[36] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6984" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2783:2736] = mn_mask_uv_lo[37] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6985" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1439:1392] = mn_mask_uv_lo[38] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6986" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2879:2832] = mn_mask_uv_lo[39] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6987" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1487:1440] = mn_mask_y_d1[20] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6988" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[2975:2928] = mn_mask_y_d1[21] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6989" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_16b_myuv[1535:1488] = mn_mask_uv_lo[40] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6990" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_8b_myuv[3071:3024] = mn_mask_uv_lo[41] ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:6991" *) 48'b000000000000000000000000000000000000000000000000 : { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign _0396_ = pk_rsp_cur_layer_end ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7293" *) sg2pack_entry_end : sg2pack_entry_mid;
  assign pk_rsp_data_entries = pk_rsp_cur_1st_height ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7293" *) sg2pack_entry_st : _0396_;
  assign _0397_ = pk_rsp_cur_layer_end ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7304" *) sg2pack_sub_h_end : sg2pack_sub_h_mid;
  assign pk_rsp_data_slices = pk_rsp_cur_1st_height ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7304" *) sg2pack_sub_h_st : _0397_;
  assign pk_rsp_wr_base_inc = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7313" *) { 1'b0, status2dma_wr_idx } : _0090_;
  assign pk_rsp_wr_base_w = is_base_wrap ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7334" *) { pk_rsp_wr_base_wrap, pk_rsp_wr_base_inc[7:0] } : pk_rsp_wr_base_inc[11:0];
  assign pk_rsp_wr_h_offset_w = _0371_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7508" *) 12'b000000000000 : _0091_;
  assign _0398_ = pixel_data_expand ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7680" *) { pk_rsp_wr_size_ori[1:0], 1'b0 } : pk_rsp_wr_size_ori;
  assign pk_rsp_wr_w_add = pixel_data_shrink ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7680" *) { 1'b0, pk_rsp_wr_size_ori[2:1] } : _0398_;
  assign _0150_[13:0] = _0148_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7694" *) pk_rsp_wr_w_offset_ori : _0092_;
  assign pk_rsp_wr_w_offset_w = _0372_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7694" *) 14'b00000000000000 : _0150_[13:0];
  assign pk_rsp_wr_addr = is_addr_wrap ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:7993" *) { pk_rsp_wr_addr_wrap, pk_rsp_wr_addr_inc[7:0] } : pk_rsp_wr_addr_inc[11:0];
  assign _0399_ = _0149_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8424" *) 1'b1 : pack_is_done;
  assign pack_is_done_w = is_first_running ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_pack.v:8424" *) 1'b0 : _0399_;
  assign _0150_[14] = 1'bx;
  assign dat_16b_yuv = { dat_l1_hi[511:480], pk_rsp_planar0_c0_d1[511:496], dat_l1_hi[479:448], pk_rsp_planar0_c0_d1[495:480], dat_l1_hi[447:416], pk_rsp_planar0_c0_d1[479:464], dat_l1_hi[415:384], pk_rsp_planar0_c0_d1[463:448], dat_l1_hi[383:352], pk_rsp_planar0_c0_d1[447:432], dat_l1_hi[351:320], pk_rsp_planar0_c0_d1[431:416], dat_l1_hi[319:288], pk_rsp_planar0_c0_d1[415:400], dat_l1_hi[287:256], pk_rsp_planar0_c0_d1[399:384], dat_l1_hi[255:224], pk_rsp_planar0_c0_d1[383:368], dat_l1_hi[223:192], pk_rsp_planar0_c0_d1[367:352], dat_l1_hi[191:160], pk_rsp_planar0_c0_d1[351:336], dat_l1_hi[159:128], pk_rsp_planar0_c0_d1[335:320], dat_l1_hi[127:96], pk_rsp_planar0_c0_d1[319:304], dat_l1_hi[95:64], pk_rsp_planar0_c0_d1[303:288], dat_l1_hi[63:32], pk_rsp_planar0_c0_d1[287:272], dat_l1_hi[31:0], pk_rsp_planar0_c0_d1[271:256], dat_l1_lo[511:480], pk_rsp_planar0_c0_d1[255:240], dat_l1_lo[479:448], pk_rsp_planar0_c0_d1[239:224], dat_l1_lo[447:416], pk_rsp_planar0_c0_d1[223:208], dat_l1_lo[415:384], pk_rsp_planar0_c0_d1[207:192], dat_l1_lo[383:352], pk_rsp_planar0_c0_d1[191:176], dat_l1_lo[351:320], pk_rsp_planar0_c0_d1[175:160], dat_l1_lo[319:288], pk_rsp_planar0_c0_d1[159:144], dat_l1_lo[287:256], pk_rsp_planar0_c0_d1[143:128], dat_l1_lo[255:224], pk_rsp_planar0_c0_d1[127:112], dat_l1_lo[223:192], pk_rsp_planar0_c0_d1[111:96], dat_l1_lo[191:160], pk_rsp_planar0_c0_d1[95:80], dat_l1_lo[159:128], pk_rsp_planar0_c0_d1[79:64], dat_l1_lo[127:96], pk_rsp_planar0_c0_d1[63:48], dat_l1_lo[95:64], pk_rsp_planar0_c0_d1[47:32], dat_l1_lo[63:32], pk_rsp_planar0_c0_d1[31:16], dat_l1_lo[31:0], pk_rsp_planar0_c0_d1[15:0] };
  assign dat_8b_yuv = { dat_l1_hi[511:496], pk_rsp_planar0_c0_d1[511:504], dat_l1_hi[495:480], pk_rsp_planar0_c0_d1[503:496], dat_l1_hi[479:464], pk_rsp_planar0_c0_d1[495:488], dat_l1_hi[463:448], pk_rsp_planar0_c0_d1[487:480], dat_l1_hi[447:432], pk_rsp_planar0_c0_d1[479:472], dat_l1_hi[431:416], pk_rsp_planar0_c0_d1[471:464], dat_l1_hi[415:400], pk_rsp_planar0_c0_d1[463:456], dat_l1_hi[399:384], pk_rsp_planar0_c0_d1[455:448], dat_l1_hi[383:368], pk_rsp_planar0_c0_d1[447:440], dat_l1_hi[367:352], pk_rsp_planar0_c0_d1[439:432], dat_l1_hi[351:336], pk_rsp_planar0_c0_d1[431:424], dat_l1_hi[335:320], pk_rsp_planar0_c0_d1[423:416], dat_l1_hi[319:304], pk_rsp_planar0_c0_d1[415:408], dat_l1_hi[303:288], pk_rsp_planar0_c0_d1[407:400], dat_l1_hi[287:272], pk_rsp_planar0_c0_d1[399:392], dat_l1_hi[271:256], pk_rsp_planar0_c0_d1[391:384], dat_l1_hi[255:240], pk_rsp_planar0_c0_d1[383:376], dat_l1_hi[239:224], pk_rsp_planar0_c0_d1[375:368], dat_l1_hi[223:208], pk_rsp_planar0_c0_d1[367:360], dat_l1_hi[207:192], pk_rsp_planar0_c0_d1[359:352], dat_l1_hi[191:176], pk_rsp_planar0_c0_d1[351:344], dat_l1_hi[175:160], pk_rsp_planar0_c0_d1[343:336], dat_l1_hi[159:144], pk_rsp_planar0_c0_d1[335:328], dat_l1_hi[143:128], pk_rsp_planar0_c0_d1[327:320], dat_l1_hi[127:112], pk_rsp_planar0_c0_d1[319:312], dat_l1_hi[111:96], pk_rsp_planar0_c0_d1[311:304], dat_l1_hi[95:80], pk_rsp_planar0_c0_d1[303:296], dat_l1_hi[79:64], pk_rsp_planar0_c0_d1[295:288], dat_l1_hi[63:48], pk_rsp_planar0_c0_d1[287:280], dat_l1_hi[47:32], pk_rsp_planar0_c0_d1[279:272], dat_l1_hi[31:16], pk_rsp_planar0_c0_d1[271:264], dat_l1_hi[15:0], pk_rsp_planar0_c0_d1[263:256], dat_l1_lo[511:496], pk_rsp_planar0_c0_d1[255:248], dat_l1_lo[495:480], pk_rsp_planar0_c0_d1[247:240], dat_l1_lo[479:464], pk_rsp_planar0_c0_d1[239:232], dat_l1_lo[463:448], pk_rsp_planar0_c0_d1[231:224], dat_l1_lo[447:432], pk_rsp_planar0_c0_d1[223:216], dat_l1_lo[431:416], pk_rsp_planar0_c0_d1[215:208], dat_l1_lo[415:400], pk_rsp_planar0_c0_d1[207:200], dat_l1_lo[399:384], pk_rsp_planar0_c0_d1[199:192], dat_l1_lo[383:368], pk_rsp_planar0_c0_d1[191:184], dat_l1_lo[367:352], pk_rsp_planar0_c0_d1[183:176], dat_l1_lo[351:336], pk_rsp_planar0_c0_d1[175:168], dat_l1_lo[335:320], pk_rsp_planar0_c0_d1[167:160], dat_l1_lo[319:304], pk_rsp_planar0_c0_d1[159:152], dat_l1_lo[303:288], pk_rsp_planar0_c0_d1[151:144], dat_l1_lo[287:272], pk_rsp_planar0_c0_d1[143:136], dat_l1_lo[271:256], pk_rsp_planar0_c0_d1[135:128], dat_l1_lo[255:240], pk_rsp_planar0_c0_d1[127:120], dat_l1_lo[239:224], pk_rsp_planar0_c0_d1[119:112], dat_l1_lo[223:208], pk_rsp_planar0_c0_d1[111:104], dat_l1_lo[207:192], pk_rsp_planar0_c0_d1[103:96], dat_l1_lo[191:176], pk_rsp_planar0_c0_d1[95:88], dat_l1_lo[175:160], pk_rsp_planar0_c0_d1[87:80], dat_l1_lo[159:144], pk_rsp_planar0_c0_d1[79:72], dat_l1_lo[143:128], pk_rsp_planar0_c0_d1[71:64], dat_l1_lo[127:112], pk_rsp_planar0_c0_d1[63:56], dat_l1_lo[111:96], pk_rsp_planar0_c0_d1[55:48], dat_l1_lo[95:80], pk_rsp_planar0_c0_d1[47:40], dat_l1_lo[79:64], pk_rsp_planar0_c0_d1[39:32], dat_l1_lo[63:48], pk_rsp_planar0_c0_d1[31:24], dat_l1_lo[47:32], pk_rsp_planar0_c0_d1[23:16], dat_l1_lo[31:16], pk_rsp_planar0_c0_d1[15:8], dat_l1_lo[15:0], pk_rsp_planar0_c0_d1[7:0] };
  assign dat_l0 = pk_rsp_planar0_c0_d1;
  assign dat_l1 = { dat_l1_hi, dat_l1_lo };
  assign dat_yuv[1535:1520] = dat_l1_hi[511:496];
  assign data_planar0_en = rd_planar0_en;
  assign data_planar0_ori_en = is_first_running;
  assign data_planar1_en = rd_planar1_en;
  assign data_planar1_ori_en = is_first_running;
  assign data_width_mark_0 = { 9'b000000000, pad_left_d1 };
  assign img2cvt_dat_wr_addr = pk_out_addr;
  assign img2cvt_dat_wr_data = { pk_out_data_h1, pk_out_data_h0 };
  assign img2cvt_dat_wr_en = pk_out_vld;
  assign img2cvt_dat_wr_hsel = pk_out_hsel;
  assign img2cvt_dat_wr_info_pd = { pk_out_sub_h, pk_out_uint, pk_out_mean, pk_out_ext128, pk_out_ext64, 1'b0, pk_out_mask };
  assign img2cvt_dat_wr_pad_mask = { pk_out_pad_mask_h1, pk_out_pad_mask_h0 };
  assign img2cvt_mn_wr_data = { pk_mn_out_data_h1, pk_mn_out_data_h0 };
  assign img2sbuf_p0_rd_addr = rd_p0_addr_d1;
  assign img2sbuf_p0_rd_en = rd_p0_vld_d1;
  assign img2sbuf_p1_rd_addr = rd_p1_addr_d1;
  assign img2sbuf_p1_rd_en = rd_p1_vld_d1;
  assign img2status_dat_entries = pk_out_data_entries;
  assign img2status_dat_slices = { 8'b00000000, pk_out_data_slices };
  assign img2status_dat_updt = pk_out_data_updt;
  assign img_layer_end = img_pd[10];
  assign img_line_end = img_pd[9];
  assign img_p0_burst = img_pd[3:0];
  assign img_p1_burst = img_pd[8:4];
  assign is_last_sub_h = 1'b1;
  assign mask_pad = { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 };
  assign mask_zero = { rd_p1_zero_mask_d3, rd_p0_zero_mask_d3 };
  assign mn_8b_mnorm[15:0] = mn_16b_mnorm[15:0];
  assign { mn_8b_myuv[3023:2976], mn_8b_myuv[2927:2880], mn_8b_myuv[2831:2784], mn_8b_myuv[2735:2688], mn_8b_myuv[2639:2592], mn_8b_myuv[2543:2496], mn_8b_myuv[2447:2400], mn_8b_myuv[2351:2304], mn_8b_myuv[2255:2208], mn_8b_myuv[2159:2112], mn_8b_myuv[2063:2016], mn_8b_myuv[1967:1920], mn_8b_myuv[1871:1824], mn_8b_myuv[1775:1728], mn_8b_myuv[1679:1632], mn_8b_myuv[1583:1536], mn_8b_myuv[1487:1440], mn_8b_myuv[1391:1344], mn_8b_myuv[1295:1248], mn_8b_myuv[1199:1152], mn_8b_myuv[1103:1056], mn_8b_myuv[1007:960], mn_8b_myuv[911:864], mn_8b_myuv[815:768], mn_8b_myuv[719:672], mn_8b_myuv[623:576], mn_8b_myuv[527:480], mn_8b_myuv[431:384], mn_8b_myuv[335:288], mn_8b_myuv[239:192], mn_8b_myuv[143:96], mn_8b_myuv[47:0] } = mn_16b_myuv;
  assign mn_ch1 = { reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry, reg2dp_mean_ry };
  assign mn_ch3 = { reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_ch4 = { reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry, reg2dp_mean_ax, reg2dp_mean_bv, reg2dp_mean_gu, reg2dp_mean_ry };
  assign mn_mask_uv[63:0] = mn_mask_uv_lo;
  assign mn_mask_uv_1_en = pk_rsp_planar1_c1_en;
  assign mn_mask_uv_hi = mn_mask_uv[127:64];
  assign mn_mask_y = mn_mask_y_d1;
  assign mn_mask_yuv = { mn_mask_y_d1[63:62], mn_mask_uv[123:120], mn_mask_y_d1[61:60], mn_mask_uv[119:116], mn_mask_y_d1[59:58], mn_mask_uv[115:112], mn_mask_y_d1[57:56], mn_mask_uv[111:108], mn_mask_y_d1[55:54], mn_mask_uv[107:104], mn_mask_y_d1[53:52], mn_mask_uv[103:100], mn_mask_y_d1[51:50], mn_mask_uv[99:96], mn_mask_y_d1[49:48], mn_mask_uv[95:92], mn_mask_y_d1[47:46], mn_mask_uv[91:88], mn_mask_y_d1[45:44], mn_mask_uv[87:84], mn_mask_y_d1[43:42], mn_mask_uv[83:80], mn_mask_y_d1[41:40], mn_mask_uv[79:76], mn_mask_y_d1[39:38], mn_mask_uv[75:72], mn_mask_y_d1[37:36], mn_mask_uv[71:68], mn_mask_y_d1[35:34], mn_mask_uv[67:64], mn_mask_y_d1[33:32], mn_mask_uv_lo[63:60], mn_mask_y_d1[31:30], mn_mask_uv_lo[59:56], mn_mask_y_d1[29:28], mn_mask_uv_lo[55:52], mn_mask_y_d1[27:26], mn_mask_uv_lo[51:48], mn_mask_y_d1[25:24], mn_mask_uv_lo[47:44], mn_mask_y_d1[23:22], mn_mask_uv_lo[43:40], mn_mask_y_d1[21:20], mn_mask_uv_lo[39:36], mn_mask_y_d1[19:18], mn_mask_uv_lo[35:32], mn_mask_y_d1[17:16], mn_mask_uv_lo[31:28], mn_mask_y_d1[15:14], mn_mask_uv_lo[27:24], mn_mask_y_d1[13:12], mn_mask_uv_lo[23:20], mn_mask_y_d1[11:10], mn_mask_uv_lo[19:16], mn_mask_y_d1[9:8], mn_mask_uv_lo[15:12], mn_mask_y_d1[7:6], mn_mask_uv_lo[11:8], mn_mask_y_d1[5:4], mn_mask_uv_lo[7:4], mn_mask_y_d1[3:2], mn_mask_uv_lo[3:0], mn_mask_y_d1[1:0] };
  assign mon_pk_rsp_wr_cnt_w = 1'bx;
  assign mon_pk_rsp_wr_h_offset_w = 1'bx;
  assign mon_pk_rsp_wr_w_offset_w = 1'bx;
  assign pad_mask_16b_yuv = { pad_mask_l1_hi[63:60], mask_pad_planar0_c0_d1[63:62], pad_mask_l1_hi[59:56], mask_pad_planar0_c0_d1[61:60], pad_mask_l1_hi[55:52], mask_pad_planar0_c0_d1[59:58], pad_mask_l1_hi[51:48], mask_pad_planar0_c0_d1[57:56], pad_mask_l1_hi[47:44], mask_pad_planar0_c0_d1[55:54], pad_mask_l1_hi[43:40], mask_pad_planar0_c0_d1[53:52], pad_mask_l1_hi[39:36], mask_pad_planar0_c0_d1[51:50], pad_mask_l1_hi[35:32], mask_pad_planar0_c0_d1[49:48], pad_mask_l1_hi[31:28], mask_pad_planar0_c0_d1[47:46], pad_mask_l1_hi[27:24], mask_pad_planar0_c0_d1[45:44], pad_mask_l1_hi[23:20], mask_pad_planar0_c0_d1[43:42], pad_mask_l1_hi[19:16], mask_pad_planar0_c0_d1[41:40], pad_mask_l1_hi[15:12], mask_pad_planar0_c0_d1[39:38], pad_mask_l1_hi[11:8], mask_pad_planar0_c0_d1[37:36], pad_mask_l1_hi[7:4], mask_pad_planar0_c0_d1[35:34], pad_mask_l1_hi[3:0], mask_pad_planar0_c0_d1[33:32], pad_mask_l1_lo[63:60], mask_pad_planar0_c0_d1[31:30], pad_mask_l1_lo[59:56], mask_pad_planar0_c0_d1[29:28], pad_mask_l1_lo[55:52], mask_pad_planar0_c0_d1[27:26], pad_mask_l1_lo[51:48], mask_pad_planar0_c0_d1[25:24], pad_mask_l1_lo[47:44], mask_pad_planar0_c0_d1[23:22], pad_mask_l1_lo[43:40], mask_pad_planar0_c0_d1[21:20], pad_mask_l1_lo[39:36], mask_pad_planar0_c0_d1[19:18], pad_mask_l1_lo[35:32], mask_pad_planar0_c0_d1[17:16], pad_mask_l1_lo[31:28], mask_pad_planar0_c0_d1[15:14], pad_mask_l1_lo[27:24], mask_pad_planar0_c0_d1[13:12], pad_mask_l1_lo[23:20], mask_pad_planar0_c0_d1[11:10], pad_mask_l1_lo[19:16], mask_pad_planar0_c0_d1[9:8], pad_mask_l1_lo[15:12], mask_pad_planar0_c0_d1[7:6], pad_mask_l1_lo[11:8], mask_pad_planar0_c0_d1[5:4], pad_mask_l1_lo[7:4], mask_pad_planar0_c0_d1[3:2], pad_mask_l1_lo[3:0], mask_pad_planar0_c0_d1[1:0] };
  assign pad_mask_8b_yuv = { pad_mask_l1_hi[63:62], mask_pad_planar0_c0_d1[63], pad_mask_l1_hi[61:60], mask_pad_planar0_c0_d1[62], pad_mask_l1_hi[59:58], mask_pad_planar0_c0_d1[61], pad_mask_l1_hi[57:56], mask_pad_planar0_c0_d1[60], pad_mask_l1_hi[55:54], mask_pad_planar0_c0_d1[59], pad_mask_l1_hi[53:52], mask_pad_planar0_c0_d1[58], pad_mask_l1_hi[51:50], mask_pad_planar0_c0_d1[57], pad_mask_l1_hi[49:48], mask_pad_planar0_c0_d1[56], pad_mask_l1_hi[47:46], mask_pad_planar0_c0_d1[55], pad_mask_l1_hi[45:44], mask_pad_planar0_c0_d1[54], pad_mask_l1_hi[43:42], mask_pad_planar0_c0_d1[53], pad_mask_l1_hi[41:40], mask_pad_planar0_c0_d1[52], pad_mask_l1_hi[39:38], mask_pad_planar0_c0_d1[51], pad_mask_l1_hi[37:36], mask_pad_planar0_c0_d1[50], pad_mask_l1_hi[35:34], mask_pad_planar0_c0_d1[49], pad_mask_l1_hi[33:32], mask_pad_planar0_c0_d1[48], pad_mask_l1_hi[31:30], mask_pad_planar0_c0_d1[47], pad_mask_l1_hi[29:28], mask_pad_planar0_c0_d1[46], pad_mask_l1_hi[27:26], mask_pad_planar0_c0_d1[45], pad_mask_l1_hi[25:24], mask_pad_planar0_c0_d1[44], pad_mask_l1_hi[23:22], mask_pad_planar0_c0_d1[43], pad_mask_l1_hi[21:20], mask_pad_planar0_c0_d1[42], pad_mask_l1_hi[19:18], mask_pad_planar0_c0_d1[41], pad_mask_l1_hi[17:16], mask_pad_planar0_c0_d1[40], pad_mask_l1_hi[15:14], mask_pad_planar0_c0_d1[39], pad_mask_l1_hi[13:12], mask_pad_planar0_c0_d1[38], pad_mask_l1_hi[11:10], mask_pad_planar0_c0_d1[37], pad_mask_l1_hi[9:8], mask_pad_planar0_c0_d1[36], pad_mask_l1_hi[7:6], mask_pad_planar0_c0_d1[35], pad_mask_l1_hi[5:4], mask_pad_planar0_c0_d1[34], pad_mask_l1_hi[3:2], mask_pad_planar0_c0_d1[33], pad_mask_l1_hi[1:0], mask_pad_planar0_c0_d1[32], pad_mask_l1_lo[63:62], mask_pad_planar0_c0_d1[31], pad_mask_l1_lo[61:60], mask_pad_planar0_c0_d1[30], pad_mask_l1_lo[59:58], mask_pad_planar0_c0_d1[29], pad_mask_l1_lo[57:56], mask_pad_planar0_c0_d1[28], pad_mask_l1_lo[55:54], mask_pad_planar0_c0_d1[27], pad_mask_l1_lo[53:52], mask_pad_planar0_c0_d1[26], pad_mask_l1_lo[51:50], mask_pad_planar0_c0_d1[25], pad_mask_l1_lo[49:48], mask_pad_planar0_c0_d1[24], pad_mask_l1_lo[47:46], mask_pad_planar0_c0_d1[23], pad_mask_l1_lo[45:44], mask_pad_planar0_c0_d1[22], pad_mask_l1_lo[43:42], mask_pad_planar0_c0_d1[21], pad_mask_l1_lo[41:40], mask_pad_planar0_c0_d1[20], pad_mask_l1_lo[39:38], mask_pad_planar0_c0_d1[19], pad_mask_l1_lo[37:36], mask_pad_planar0_c0_d1[18], pad_mask_l1_lo[35:34], mask_pad_planar0_c0_d1[17], pad_mask_l1_lo[33:32], mask_pad_planar0_c0_d1[16], pad_mask_l1_lo[31:30], mask_pad_planar0_c0_d1[15], pad_mask_l1_lo[29:28], mask_pad_planar0_c0_d1[14], pad_mask_l1_lo[27:26], mask_pad_planar0_c0_d1[13], pad_mask_l1_lo[25:24], mask_pad_planar0_c0_d1[12], pad_mask_l1_lo[23:22], mask_pad_planar0_c0_d1[11], pad_mask_l1_lo[21:20], mask_pad_planar0_c0_d1[10], pad_mask_l1_lo[19:18], mask_pad_planar0_c0_d1[9], pad_mask_l1_lo[17:16], mask_pad_planar0_c0_d1[8], pad_mask_l1_lo[15:14], mask_pad_planar0_c0_d1[7], pad_mask_l1_lo[13:12], mask_pad_planar0_c0_d1[6], pad_mask_l1_lo[11:10], mask_pad_planar0_c0_d1[5], pad_mask_l1_lo[9:8], mask_pad_planar0_c0_d1[4], pad_mask_l1_lo[7:6], mask_pad_planar0_c0_d1[3], pad_mask_l1_lo[5:4], mask_pad_planar0_c0_d1[2], pad_mask_l1_lo[3:2], mask_pad_planar0_c0_d1[1], pad_mask_l1_lo[1:0], mask_pad_planar0_c0_d1[0] };
  assign pad_mask_l0 = mask_pad_planar0_c0_d1;
  assign pad_mask_l1 = { pad_mask_l1_hi, pad_mask_l1_lo };
  assign pad_mask_yuv[191:190] = pad_mask_l1_hi[63:62];
  assign pk_mn_out_data = { pk_mn_out_data_h1, pk_mn_out_data_h0 };
  assign pk_out_data = { pk_out_data_h1, pk_out_data_h0 };
  assign pk_out_info_pd = { pk_out_sub_h, pk_out_uint, pk_out_mean, pk_out_ext128, pk_out_ext64, 1'b0, pk_out_mask };
  assign pk_out_interleave = 1'b0;
  assign pk_out_pad_mask = { pk_out_pad_mask_h1, pk_out_pad_mask_h0 };
  assign pk_rsp_1st_height = rd_1st_height_d3;
  assign pk_rsp_cur_vld = pk_rsp_wr_vld;
  assign pk_rsp_dat_ergb = { img2sbuf_p1_rd_data[255:254], 14'b00000000000000, img2sbuf_p1_rd_data[253:244], 6'b000000, img2sbuf_p1_rd_data[243:234], 6'b000000, img2sbuf_p1_rd_data[233:224], 6'b000000, img2sbuf_p1_rd_data[223:222], 14'b00000000000000, img2sbuf_p1_rd_data[221:212], 6'b000000, img2sbuf_p1_rd_data[211:202], 6'b000000, img2sbuf_p1_rd_data[201:192], 6'b000000, img2sbuf_p1_rd_data[191:190], 14'b00000000000000, img2sbuf_p1_rd_data[189:180], 6'b000000, img2sbuf_p1_rd_data[179:170], 6'b000000, img2sbuf_p1_rd_data[169:160], 6'b000000, img2sbuf_p1_rd_data[159:158], 14'b00000000000000, img2sbuf_p1_rd_data[157:148], 6'b000000, img2sbuf_p1_rd_data[147:138], 6'b000000, img2sbuf_p1_rd_data[137:128], 6'b000000, img2sbuf_p1_rd_data[127:126], 14'b00000000000000, img2sbuf_p1_rd_data[125:116], 6'b000000, img2sbuf_p1_rd_data[115:106], 6'b000000, img2sbuf_p1_rd_data[105:96], 6'b000000, img2sbuf_p1_rd_data[95:94], 14'b00000000000000, img2sbuf_p1_rd_data[93:84], 6'b000000, img2sbuf_p1_rd_data[83:74], 6'b000000, img2sbuf_p1_rd_data[73:64], 6'b000000, img2sbuf_p1_rd_data[63:62], 14'b00000000000000, img2sbuf_p1_rd_data[61:52], 6'b000000, img2sbuf_p1_rd_data[51:42], 6'b000000, img2sbuf_p1_rd_data[41:32], 6'b000000, img2sbuf_p1_rd_data[31:30], 14'b00000000000000, img2sbuf_p1_rd_data[29:20], 6'b000000, img2sbuf_p1_rd_data[19:10], 6'b000000, img2sbuf_p1_rd_data[9:0], 6'b000000, img2sbuf_p0_rd_data[255:254], 14'b00000000000000, img2sbuf_p0_rd_data[253:244], 6'b000000, img2sbuf_p0_rd_data[243:234], 6'b000000, img2sbuf_p0_rd_data[233:224], 6'b000000, img2sbuf_p0_rd_data[223:222], 14'b00000000000000, img2sbuf_p0_rd_data[221:212], 6'b000000, img2sbuf_p0_rd_data[211:202], 6'b000000, img2sbuf_p0_rd_data[201:192], 6'b000000, img2sbuf_p0_rd_data[191:190], 14'b00000000000000, img2sbuf_p0_rd_data[189:180], 6'b000000, img2sbuf_p0_rd_data[179:170], 6'b000000, img2sbuf_p0_rd_data[169:160], 6'b000000, img2sbuf_p0_rd_data[159:158], 14'b00000000000000, img2sbuf_p0_rd_data[157:148], 6'b000000, img2sbuf_p0_rd_data[147:138], 6'b000000, img2sbuf_p0_rd_data[137:128], 6'b000000, img2sbuf_p0_rd_data[127:126], 14'b00000000000000, img2sbuf_p0_rd_data[125:116], 6'b000000, img2sbuf_p0_rd_data[115:106], 6'b000000, img2sbuf_p0_rd_data[105:96], 6'b000000, img2sbuf_p0_rd_data[95:94], 14'b00000000000000, img2sbuf_p0_rd_data[93:84], 6'b000000, img2sbuf_p0_rd_data[83:74], 6'b000000, img2sbuf_p0_rd_data[73:64], 6'b000000, img2sbuf_p0_rd_data[63:62], 14'b00000000000000, img2sbuf_p0_rd_data[61:52], 6'b000000, img2sbuf_p0_rd_data[51:42], 6'b000000, img2sbuf_p0_rd_data[41:32], 6'b000000, img2sbuf_p0_rd_data[31:30], 14'b00000000000000, img2sbuf_p0_rd_data[29:20], 6'b000000, img2sbuf_p0_rd_data[19:10], 6'b000000, img2sbuf_p0_rd_data[9:0], 6'b000000 };
  assign pk_rsp_dat_mergb[1023:512] = pk_rsp_data_h1;
  assign pk_rsp_dat_normal = { img2sbuf_p1_rd_data, img2sbuf_p0_rd_data };
  assign pk_rsp_data_h0_en = pk_rsp_wr_vld;
  assign pk_rsp_layer_end = rd_layer_end_d3;
  assign pk_rsp_loop_end = rd_loop_end_d3;
  assign pk_rsp_mn_data_h0_en = pk_rsp_wr_vld;
  assign pk_rsp_one_line_end = rd_one_line_end_d3;
  assign pk_rsp_out_sel[0] = pixel_packed_10b;
  assign pk_rsp_p0_data = img2sbuf_p0_rd_data;
  assign pk_rsp_p0_pad_mask = rd_p0_pad_mask_d3;
  assign pk_rsp_p0_zero_mask = rd_p0_zero_mask_d3;
  assign pk_rsp_p1_data = img2sbuf_p1_rd_data;
  assign pk_rsp_p1_pad_mask = rd_p1_pad_mask_d3;
  assign pk_rsp_p1_zero_mask = rd_p1_zero_mask_d3;
  assign pk_rsp_pad_mask_ergb = { rd_p1_pad_mask_d3[31], rd_p1_pad_mask_d3[31:30], rd_p1_pad_mask_d3[30:29], rd_p1_pad_mask_d3[29:28], rd_p1_pad_mask_d3[28:27], rd_p1_pad_mask_d3[27:26], rd_p1_pad_mask_d3[26:25], rd_p1_pad_mask_d3[25:24], rd_p1_pad_mask_d3[24:23], rd_p1_pad_mask_d3[23:22], rd_p1_pad_mask_d3[22:21], rd_p1_pad_mask_d3[21:20], rd_p1_pad_mask_d3[20:19], rd_p1_pad_mask_d3[19:18], rd_p1_pad_mask_d3[18:17], rd_p1_pad_mask_d3[17:16], rd_p1_pad_mask_d3[16:15], rd_p1_pad_mask_d3[15:14], rd_p1_pad_mask_d3[14:13], rd_p1_pad_mask_d3[13:12], rd_p1_pad_mask_d3[12:11], rd_p1_pad_mask_d3[11:10], rd_p1_pad_mask_d3[10:9], rd_p1_pad_mask_d3[9:8], rd_p1_pad_mask_d3[8:7], rd_p1_pad_mask_d3[7:6], rd_p1_pad_mask_d3[6:5], rd_p1_pad_mask_d3[5:4], rd_p1_pad_mask_d3[4:3], rd_p1_pad_mask_d3[3:2], rd_p1_pad_mask_d3[2:1], rd_p1_pad_mask_d3[1:0], rd_p1_pad_mask_d3[0], rd_p0_pad_mask_d3[31], rd_p0_pad_mask_d3[31:30], rd_p0_pad_mask_d3[30:29], rd_p0_pad_mask_d3[29:28], rd_p0_pad_mask_d3[28:27], rd_p0_pad_mask_d3[27:26], rd_p0_pad_mask_d3[26:25], rd_p0_pad_mask_d3[25:24], rd_p0_pad_mask_d3[24:23], rd_p0_pad_mask_d3[23:22], rd_p0_pad_mask_d3[22:21], rd_p0_pad_mask_d3[21:20], rd_p0_pad_mask_d3[20:19], rd_p0_pad_mask_d3[19:18], rd_p0_pad_mask_d3[18:17], rd_p0_pad_mask_d3[17:16], rd_p0_pad_mask_d3[16:15], rd_p0_pad_mask_d3[15:14], rd_p0_pad_mask_d3[14:13], rd_p0_pad_mask_d3[13:12], rd_p0_pad_mask_d3[12:11], rd_p0_pad_mask_d3[11:10], rd_p0_pad_mask_d3[10:9], rd_p0_pad_mask_d3[9:8], rd_p0_pad_mask_d3[8:7], rd_p0_pad_mask_d3[7:6], rd_p0_pad_mask_d3[6:5], rd_p0_pad_mask_d3[5:4], rd_p0_pad_mask_d3[4:3], rd_p0_pad_mask_d3[3:2], rd_p0_pad_mask_d3[2:1], rd_p0_pad_mask_d3[1:0], rd_p0_pad_mask_d3[0] };
  assign pk_rsp_pad_mask_norm = { rd_p1_pad_mask_d3, rd_p0_pad_mask_d3 };
  assign pk_rsp_planar = rd_planar_d3;
  assign pk_rsp_planar0_c0_en = mn_mask_y_en;
  assign pk_rsp_planar1_c0_en = mn_mask_uv_0_en;
  assign pk_rsp_sub_h = rd_sub_h_d3;
  assign pk_rsp_sub_h_end = rd_sub_h_end_d3;
  assign pk_rsp_vld = rd_vld_d3;
  assign pk_rsp_wr_entries = pk_rsp_data_entries;
  assign pk_rsp_wr_slices = pk_rsp_data_slices;
  assign pk_rsp_wr_sub_addr = pk_rsp_wr_w_offset[1:0];
  assign pk_rsp_wr_w_offset_ori_en = is_first_running;
  assign rd_planar0_ori_en = is_first_running;
  assign rd_planar1_ori_en = is_first_running;
  assign rd_sub_h_cnt = 3'b000;
  assign rd_sub_h_end = rd_loop_end;
  assign rdat = { img2sbuf_p1_rd_data, img2sbuf_p0_rd_data };
  assign z14 = 14'b00000000000000;
  assign z6 = 6'b000000;
endmodule
