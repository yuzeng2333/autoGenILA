module CDP_ICVT_chn_data_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:241" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:242" *)
  output outsig;
  assign outsig = in_0;
endmodule
