module NV_NVDLA_cbuf(nvdla_core_clk, nvdla_core_rstn, cdma2buf_dat_wr_addr, cdma2buf_dat_wr_data, cdma2buf_dat_wr_en, cdma2buf_dat_wr_hsel, cdma2buf_wt_wr_addr, cdma2buf_wt_wr_data, cdma2buf_wt_wr_en, cdma2buf_wt_wr_hsel, pwrbus_ram_pd, sc2buf_dat_rd_addr, sc2buf_dat_rd_en, sc2buf_wmb_rd_addr, sc2buf_wmb_rd_en, sc2buf_wt_rd_addr, sc2buf_wt_rd_en, sc2buf_dat_rd_data, sc2buf_dat_rd_valid, sc2buf_wmb_rd_data, sc2buf_wmb_rd_valid, sc2buf_wt_rd_data, sc2buf_wt_rd_valid);
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5719" *)
  wire [511:0] _0000_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5738" *)
  wire [511:0] _0001_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5647" *)
  wire [511:0] _0002_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5637" *)
  wire [511:0] _0003_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5871" *)
  wire [511:0] _0004_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5876" *)
  wire [511:0] _0005_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1565" *)
  wire [7:0] _0006_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1595" *)
  wire [511:0] _0007_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1585" *)
  wire [511:0] _0008_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5757" *)
  wire [511:0] _0009_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5776" *)
  wire [511:0] _0010_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5667" *)
  wire [511:0] _0011_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5657" *)
  wire [511:0] _0012_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5881" *)
  wire [511:0] _0013_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5886" *)
  wire [511:0] _0014_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1575" *)
  wire [7:0] _0015_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1615" *)
  wire [511:0] _0016_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1605" *)
  wire [511:0] _0017_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5795" *)
  wire [511:0] _0018_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5814" *)
  wire [511:0] _0019_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5687" *)
  wire [511:0] _0020_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5677" *)
  wire [511:0] _0021_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5891" *)
  wire [511:0] _0022_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5896" *)
  wire [511:0] _0023_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4494" *)
  wire [7:0] _0024_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4504" *)
  wire [7:0] _0025_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4694" *)
  wire [7:0] _0026_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4704" *)
  wire [7:0] _0027_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4714" *)
  wire [7:0] _0028_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4724" *)
  wire [7:0] _0029_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4734" *)
  wire [7:0] _0030_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4744" *)
  wire [7:0] _0031_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4754" *)
  wire [7:0] _0032_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4764" *)
  wire [7:0] _0033_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4774" *)
  wire [7:0] _0034_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4784" *)
  wire [7:0] _0035_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4794" *)
  wire [7:0] _0036_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4804" *)
  wire [7:0] _0037_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4514" *)
  wire [7:0] _0038_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4524" *)
  wire [7:0] _0039_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4534" *)
  wire [7:0] _0040_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4544" *)
  wire [7:0] _0041_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4554" *)
  wire [7:0] _0042_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4564" *)
  wire [7:0] _0043_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4574" *)
  wire [7:0] _0044_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4584" *)
  wire [7:0] _0045_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4594" *)
  wire [7:0] _0046_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4604" *)
  wire [7:0] _0047_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4614" *)
  wire [7:0] _0048_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4624" *)
  wire [7:0] _0049_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4634" *)
  wire [7:0] _0050_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4644" *)
  wire [7:0] _0051_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4654" *)
  wire [7:0] _0052_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4664" *)
  wire [7:0] _0053_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4674" *)
  wire [7:0] _0054_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4684" *)
  wire [7:0] _0055_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5075" *)
  wire [511:0] _0056_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5085" *)
  wire [511:0] _0057_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5275" *)
  wire [511:0] _0058_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5285" *)
  wire [511:0] _0059_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5295" *)
  wire [511:0] _0060_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5305" *)
  wire [511:0] _0061_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5315" *)
  wire [511:0] _0062_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5325" *)
  wire [511:0] _0063_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5335" *)
  wire [511:0] _0064_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5345" *)
  wire [511:0] _0065_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5355" *)
  wire [511:0] _0066_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5365" *)
  wire [511:0] _0067_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5375" *)
  wire [511:0] _0068_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5385" *)
  wire [511:0] _0069_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5095" *)
  wire [511:0] _0070_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5105" *)
  wire [511:0] _0071_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5115" *)
  wire [511:0] _0072_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5125" *)
  wire [511:0] _0073_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5135" *)
  wire [511:0] _0074_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5145" *)
  wire [511:0] _0075_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5155" *)
  wire [511:0] _0076_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5165" *)
  wire [511:0] _0077_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5175" *)
  wire [511:0] _0078_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5185" *)
  wire [511:0] _0079_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5195" *)
  wire [511:0] _0080_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5205" *)
  wire [511:0] _0081_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5215" *)
  wire [511:0] _0082_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5225" *)
  wire [511:0] _0083_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5235" *)
  wire [511:0] _0084_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5245" *)
  wire [511:0] _0085_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5255" *)
  wire [511:0] _0086_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5265" *)
  wire [511:0] _0087_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2311" *)
  wire [7:0] _0088_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2321" *)
  wire [7:0] _0089_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2511" *)
  wire [7:0] _0090_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2521" *)
  wire [7:0] _0091_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2531" *)
  wire [7:0] _0092_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2541" *)
  wire [7:0] _0093_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2551" *)
  wire [7:0] _0094_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2561" *)
  wire [7:0] _0095_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2571" *)
  wire [7:0] _0096_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2581" *)
  wire [7:0] _0097_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2591" *)
  wire [7:0] _0098_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2601" *)
  wire [7:0] _0099_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2611" *)
  wire [7:0] _0100_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2621" *)
  wire [7:0] _0101_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2331" *)
  wire [7:0] _0102_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2341" *)
  wire [7:0] _0103_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2351" *)
  wire [7:0] _0104_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2361" *)
  wire [7:0] _0105_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2371" *)
  wire [7:0] _0106_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2381" *)
  wire [7:0] _0107_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2391" *)
  wire [7:0] _0108_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2401" *)
  wire [7:0] _0109_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2411" *)
  wire [7:0] _0110_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2421" *)
  wire [7:0] _0111_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2431" *)
  wire [7:0] _0112_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2441" *)
  wire [7:0] _0113_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2451" *)
  wire [7:0] _0114_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2461" *)
  wire [7:0] _0115_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2471" *)
  wire [7:0] _0116_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2481" *)
  wire [7:0] _0117_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2491" *)
  wire [7:0] _0118_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2501" *)
  wire [7:0] _0119_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2631" *)
  wire [511:0] _0120_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2641" *)
  wire [511:0] _0121_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2831" *)
  wire [511:0] _0122_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2841" *)
  wire [511:0] _0123_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2851" *)
  wire [511:0] _0124_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2861" *)
  wire [511:0] _0125_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2871" *)
  wire [511:0] _0126_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2881" *)
  wire [511:0] _0127_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2891" *)
  wire [511:0] _0128_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2901" *)
  wire [511:0] _0129_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2911" *)
  wire [511:0] _0130_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2921" *)
  wire [511:0] _0131_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2931" *)
  wire [511:0] _0132_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2941" *)
  wire [511:0] _0133_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2651" *)
  wire [511:0] _0134_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2661" *)
  wire [511:0] _0135_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2671" *)
  wire [511:0] _0136_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2681" *)
  wire [511:0] _0137_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2691" *)
  wire [511:0] _0138_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2701" *)
  wire [511:0] _0139_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2711" *)
  wire [511:0] _0140_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2721" *)
  wire [511:0] _0141_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2731" *)
  wire [511:0] _0142_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2741" *)
  wire [511:0] _0143_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2751" *)
  wire [511:0] _0144_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2761" *)
  wire [511:0] _0145_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2771" *)
  wire [511:0] _0146_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2781" *)
  wire [511:0] _0147_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2791" *)
  wire [511:0] _0148_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2801" *)
  wire [511:0] _0149_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2811" *)
  wire [511:0] _0150_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2821" *)
  wire [511:0] _0151_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1481" *)
  wire _0152_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1488" *)
  wire _0153_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1495" *)
  wire _0154_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1502" *)
  wire _0155_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1509" *)
  wire _0156_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1516" *)
  wire _0157_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1523" *)
  wire _0158_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1530" *)
  wire _0159_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1537" *)
  wire _0160_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1544" *)
  wire _0161_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1355" *)
  wire _0162_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1362" *)
  wire _0163_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1369" *)
  wire _0164_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1376" *)
  wire _0165_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1383" *)
  wire _0166_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1390" *)
  wire _0167_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1397" *)
  wire _0168_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1404" *)
  wire _0169_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1411" *)
  wire _0170_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1418" *)
  wire _0171_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1425" *)
  wire _0172_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1432" *)
  wire _0173_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1439" *)
  wire _0174_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1446" *)
  wire _0175_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1453" *)
  wire _0176_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1460" *)
  wire _0177_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1467" *)
  wire _0178_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1474" *)
  wire _0179_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1712" *)
  wire [7:0] _0180_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1713" *)
  wire [7:0] _0181_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1714" *)
  wire [511:0] _0182_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1715" *)
  wire [511:0] _0183_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1725" *)
  wire [7:0] _0184_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1726" *)
  wire [7:0] _0185_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1727" *)
  wire [511:0] _0186_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1728" *)
  wire [511:0] _0187_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1738" *)
  wire [7:0] _0188_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1739" *)
  wire [7:0] _0189_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1740" *)
  wire [511:0] _0190_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1741" *)
  wire [511:0] _0191_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1751" *)
  wire [7:0] _0192_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1752" *)
  wire [7:0] _0193_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1753" *)
  wire [511:0] _0194_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1754" *)
  wire [511:0] _0195_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1764" *)
  wire [7:0] _0196_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1765" *)
  wire [7:0] _0197_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1766" *)
  wire [511:0] _0198_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1767" *)
  wire [511:0] _0199_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1777" *)
  wire [7:0] _0200_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1778" *)
  wire [7:0] _0201_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1779" *)
  wire [511:0] _0202_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1780" *)
  wire [511:0] _0203_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1790" *)
  wire [7:0] _0204_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1791" *)
  wire [7:0] _0205_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1792" *)
  wire [511:0] _0206_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1793" *)
  wire [511:0] _0207_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1803" *)
  wire [7:0] _0208_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1804" *)
  wire [7:0] _0209_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1805" *)
  wire [511:0] _0210_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1806" *)
  wire [511:0] _0211_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1816" *)
  wire [7:0] _0212_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1817" *)
  wire [7:0] _0213_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1818" *)
  wire [511:0] _0214_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1819" *)
  wire [511:0] _0215_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1829" *)
  wire [7:0] _0216_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1830" *)
  wire [7:0] _0217_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1831" *)
  wire [511:0] _0218_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1832" *)
  wire [511:0] _0219_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1842" *)
  wire [7:0] _0220_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1843" *)
  wire [7:0] _0221_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1844" *)
  wire [511:0] _0222_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1845" *)
  wire [511:0] _0223_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1855" *)
  wire [7:0] _0224_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1856" *)
  wire [7:0] _0225_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1857" *)
  wire [511:0] _0226_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1858" *)
  wire [511:0] _0227_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1868" *)
  wire [7:0] _0228_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1869" *)
  wire [7:0] _0229_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1870" *)
  wire [511:0] _0230_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1871" *)
  wire [511:0] _0231_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1881" *)
  wire [7:0] _0232_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1882" *)
  wire [7:0] _0233_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1883" *)
  wire [511:0] _0234_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1884" *)
  wire [511:0] _0235_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1894" *)
  wire [7:0] _0236_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1895" *)
  wire [7:0] _0237_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1896" *)
  wire [511:0] _0238_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1897" *)
  wire [511:0] _0239_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1907" *)
  wire [7:0] _0240_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1908" *)
  wire [7:0] _0241_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1909" *)
  wire [511:0] _0242_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1910" *)
  wire [511:0] _0243_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1920" *)
  wire [7:0] _0244_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1921" *)
  wire [7:0] _0245_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1922" *)
  wire [511:0] _0246_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1923" *)
  wire [511:0] _0247_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1933" *)
  wire [7:0] _0248_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1934" *)
  wire [7:0] _0249_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1935" *)
  wire [511:0] _0250_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1936" *)
  wire [511:0] _0251_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1946" *)
  wire [7:0] _0252_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1947" *)
  wire [7:0] _0253_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1948" *)
  wire [511:0] _0254_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1949" *)
  wire [511:0] _0255_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1959" *)
  wire [7:0] _0256_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1960" *)
  wire [7:0] _0257_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1961" *)
  wire [511:0] _0258_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1962" *)
  wire [511:0] _0259_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1972" *)
  wire [7:0] _0260_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1973" *)
  wire [7:0] _0261_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1974" *)
  wire [511:0] _0262_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1975" *)
  wire [511:0] _0263_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1985" *)
  wire [7:0] _0264_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1986" *)
  wire [7:0] _0265_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1987" *)
  wire [511:0] _0266_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1988" *)
  wire [511:0] _0267_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1998" *)
  wire [7:0] _0268_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1999" *)
  wire [7:0] _0269_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2000" *)
  wire [511:0] _0270_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2001" *)
  wire [511:0] _0271_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2011" *)
  wire [7:0] _0272_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2012" *)
  wire [7:0] _0273_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2013" *)
  wire [511:0] _0274_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2014" *)
  wire [511:0] _0275_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2024" *)
  wire [7:0] _0276_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2025" *)
  wire [7:0] _0277_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2026" *)
  wire [511:0] _0278_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2027" *)
  wire [511:0] _0279_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2037" *)
  wire [7:0] _0280_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2038" *)
  wire [7:0] _0281_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2039" *)
  wire [511:0] _0282_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2040" *)
  wire [511:0] _0283_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2050" *)
  wire [7:0] _0284_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2051" *)
  wire [7:0] _0285_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2052" *)
  wire [511:0] _0286_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2053" *)
  wire [511:0] _0287_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2063" *)
  wire [7:0] _0288_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2064" *)
  wire [7:0] _0289_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2065" *)
  wire [511:0] _0290_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2066" *)
  wire [511:0] _0291_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3926" *)
  wire [7:0] _0292_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3927" *)
  wire [7:0] _0293_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3944" *)
  wire [7:0] _0294_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3945" *)
  wire [7:0] _0295_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3962" *)
  wire [7:0] _0296_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3963" *)
  wire [7:0] _0297_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3980" *)
  wire [7:0] _0298_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3981" *)
  wire [7:0] _0299_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3998" *)
  wire [7:0] _0300_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3999" *)
  wire [7:0] _0301_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4016" *)
  wire [7:0] _0302_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4017" *)
  wire [7:0] _0303_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4034" *)
  wire [7:0] _0304_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4035" *)
  wire [7:0] _0305_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4052" *)
  wire [7:0] _0306_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4053" *)
  wire [7:0] _0307_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4070" *)
  wire [7:0] _0308_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4071" *)
  wire [7:0] _0309_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4088" *)
  wire [7:0] _0310_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4089" *)
  wire [7:0] _0311_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4106" *)
  wire [7:0] _0312_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4107" *)
  wire [7:0] _0313_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4124" *)
  wire [7:0] _0314_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4125" *)
  wire [7:0] _0315_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4142" *)
  wire [7:0] _0316_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4143" *)
  wire [7:0] _0317_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4160" *)
  wire [7:0] _0318_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4161" *)
  wire [7:0] _0319_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4178" *)
  wire [7:0] _0320_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4179" *)
  wire [7:0] _0321_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5525" *)
  wire [1023:0] _0322_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5526" *)
  wire [1023:0] _0323_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5527" *)
  wire [1023:0] _0324_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5528" *)
  wire [1023:0] _0325_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5529" *)
  wire [1023:0] _0326_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5530" *)
  wire [1023:0] _0327_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5531" *)
  wire [1023:0] _0328_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5532" *)
  wire [1023:0] _0329_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5533" *)
  wire [1023:0] _0330_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5534" *)
  wire [1023:0] _0331_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5535" *)
  wire [1023:0] _0332_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5536" *)
  wire [1023:0] _0333_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5537" *)
  wire [1023:0] _0334_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5538" *)
  wire [1023:0] _0335_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5539" *)
  wire [1023:0] _0336_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5603" *)
  wire [1023:0] _0337_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5604" *)
  wire [1023:0] _0338_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5605" *)
  wire [1023:0] _0339_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5606" *)
  wire [1023:0] _0340_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5607" *)
  wire [1023:0] _0341_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5608" *)
  wire [1023:0] _0342_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5609" *)
  wire [1023:0] _0343_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5610" *)
  wire [1023:0] _0344_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5611" *)
  wire [1023:0] _0345_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5612" *)
  wire [1023:0] _0346_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5613" *)
  wire [1023:0] _0347_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5614" *)
  wire [1023:0] _0348_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5615" *)
  wire [1023:0] _0349_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5616" *)
  wire [1023:0] _0350_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5617" *)
  wire [1023:0] _0351_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1003" *)
  wire _0352_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1010" *)
  wire _0353_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1024" *)
  wire _0354_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1038" *)
  wire _0355_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1052" *)
  wire _0356_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1066" *)
  wire _0357_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1080" *)
  wire _0358_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1094" *)
  wire _0359_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1108" *)
  wire _0360_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1122" *)
  wire _0361_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1136" *)
  wire _0362_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1150" *)
  wire _0363_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1164" *)
  wire _0364_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1178" *)
  wire _0365_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1192" *)
  wire _0366_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1206" *)
  wire _0367_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1220" *)
  wire _0368_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1234" *)
  wire _0369_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1248" *)
  wire _0370_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1262" *)
  wire _0371_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3292" *)
  wire _0372_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3306" *)
  wire _0373_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3320" *)
  wire _0374_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3334" *)
  wire _0375_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3348" *)
  wire _0376_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3362" *)
  wire _0377_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3376" *)
  wire _0378_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3390" *)
  wire _0379_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3404" *)
  wire _0380_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3418" *)
  wire _0381_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3432" *)
  wire _0382_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3446" *)
  wire _0383_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3460" *)
  wire _0384_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3474" *)
  wire _0385_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3488" *)
  wire _0386_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3502" *)
  wire _0387_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3516" *)
  wire _0388_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3530" *)
  wire _0389_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3544" *)
  wire _0390_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3558" *)
  wire _0391_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3572" *)
  wire _0392_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3586" *)
  wire _0393_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3600" *)
  wire _0394_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3614" *)
  wire _0395_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3628" *)
  wire _0396_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3642" *)
  wire _0397_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3656" *)
  wire _0398_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3670" *)
  wire _0399_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3684" *)
  wire _0400_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3698" *)
  wire _0401_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:856" *)
  wire _0402_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:870" *)
  wire _0403_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:884" *)
  wire _0404_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:898" *)
  wire _0405_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:912" *)
  wire _0406_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:926" *)
  wire _0407_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:940" *)
  wire _0408_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:954" *)
  wire _0409_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:968" *)
  wire _0410_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:982" *)
  wire _0411_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:835" *)
  wire _0412_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5526" *)
  wire [1023:0] _0413_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5527" *)
  wire [1023:0] _0414_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5528" *)
  wire [1023:0] _0415_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5529" *)
  wire [1023:0] _0416_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5530" *)
  wire [1023:0] _0417_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5531" *)
  wire [1023:0] _0418_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5532" *)
  wire [1023:0] _0419_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5533" *)
  wire [1023:0] _0420_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5534" *)
  wire [1023:0] _0421_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5535" *)
  wire [1023:0] _0422_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5536" *)
  wire [1023:0] _0423_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5537" *)
  wire [1023:0] _0424_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5538" *)
  wire [1023:0] _0425_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5604" *)
  wire [1023:0] _0426_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5605" *)
  wire [1023:0] _0427_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5606" *)
  wire [1023:0] _0428_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5607" *)
  wire [1023:0] _0429_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5608" *)
  wire [1023:0] _0430_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5609" *)
  wire [1023:0] _0431_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5610" *)
  wire [1023:0] _0432_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5611" *)
  wire [1023:0] _0433_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5612" *)
  wire [1023:0] _0434_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5613" *)
  wire [1023:0] _0435_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5614" *)
  wire [1023:0] _0436_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5615" *)
  wire [1023:0] _0437_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5616" *)
  wire [1023:0] _0438_;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:61" *)
  wire [11:0] cbuf_p0_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:62" *)
  wire [3:0] cbuf_p0_rd_bank;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:63" *)
  wire [511:0] cbuf_p0_rd_c0_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:268" *)
  reg [511:0] cbuf_p0_rd_c0_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:64" *)
  wire [511:0] cbuf_p0_rd_c0_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:269" *)
  wire cbuf_p0_rd_c0_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:65" *)
  wire cbuf_p0_rd_c0_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:66" *)
  wire [511:0] cbuf_p0_rd_c1_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:270" *)
  reg [511:0] cbuf_p0_rd_c1_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:67" *)
  wire [511:0] cbuf_p0_rd_c1_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:271" *)
  wire cbuf_p0_rd_c1_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:68" *)
  wire cbuf_p0_rd_c1_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:272" *)
  reg [1023:0] cbuf_p0_rd_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:273" *)
  wire [1023:0] cbuf_p0_rd_data_d4_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:274" *)
  reg [1023:0] cbuf_p0_rd_data_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:69" *)
  wire cbuf_p0_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:70" *)
  wire cbuf_p0_rd_en_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:71" *)
  wire cbuf_p0_rd_en_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:275" *)
  reg cbuf_p0_rd_en_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:72" *)
  wire cbuf_p0_rd_sel_ram_b0c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:276" *)
  wire cbuf_p0_rd_sel_ram_b0c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:73" *)
  wire cbuf_p0_rd_sel_ram_b0c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:277" *)
  wire cbuf_p0_rd_sel_ram_b0c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:74" *)
  wire cbuf_p0_rd_sel_ram_b10c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:278" *)
  wire cbuf_p0_rd_sel_ram_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:75" *)
  wire cbuf_p0_rd_sel_ram_b10c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:279" *)
  wire cbuf_p0_rd_sel_ram_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:76" *)
  wire cbuf_p0_rd_sel_ram_b11c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:280" *)
  wire cbuf_p0_rd_sel_ram_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:77" *)
  wire cbuf_p0_rd_sel_ram_b11c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:281" *)
  wire cbuf_p0_rd_sel_ram_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:78" *)
  wire cbuf_p0_rd_sel_ram_b12c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:282" *)
  wire cbuf_p0_rd_sel_ram_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:79" *)
  wire cbuf_p0_rd_sel_ram_b12c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:283" *)
  wire cbuf_p0_rd_sel_ram_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:80" *)
  wire cbuf_p0_rd_sel_ram_b13c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:284" *)
  wire cbuf_p0_rd_sel_ram_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:81" *)
  wire cbuf_p0_rd_sel_ram_b13c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:285" *)
  wire cbuf_p0_rd_sel_ram_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:82" *)
  wire cbuf_p0_rd_sel_ram_b14c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:286" *)
  wire cbuf_p0_rd_sel_ram_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:83" *)
  wire cbuf_p0_rd_sel_ram_b14c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:287" *)
  wire cbuf_p0_rd_sel_ram_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:84" *)
  wire cbuf_p0_rd_sel_ram_b1c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:288" *)
  wire cbuf_p0_rd_sel_ram_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:85" *)
  wire cbuf_p0_rd_sel_ram_b1c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:289" *)
  wire cbuf_p0_rd_sel_ram_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:86" *)
  wire cbuf_p0_rd_sel_ram_b2c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:290" *)
  wire cbuf_p0_rd_sel_ram_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:87" *)
  wire cbuf_p0_rd_sel_ram_b2c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:291" *)
  wire cbuf_p0_rd_sel_ram_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:88" *)
  wire cbuf_p0_rd_sel_ram_b3c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:292" *)
  wire cbuf_p0_rd_sel_ram_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:89" *)
  wire cbuf_p0_rd_sel_ram_b3c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:293" *)
  wire cbuf_p0_rd_sel_ram_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:90" *)
  wire cbuf_p0_rd_sel_ram_b4c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:294" *)
  wire cbuf_p0_rd_sel_ram_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:91" *)
  wire cbuf_p0_rd_sel_ram_b4c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:295" *)
  wire cbuf_p0_rd_sel_ram_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:92" *)
  wire cbuf_p0_rd_sel_ram_b5c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:296" *)
  wire cbuf_p0_rd_sel_ram_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:93" *)
  wire cbuf_p0_rd_sel_ram_b5c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:297" *)
  wire cbuf_p0_rd_sel_ram_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:94" *)
  wire cbuf_p0_rd_sel_ram_b6c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:298" *)
  wire cbuf_p0_rd_sel_ram_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:95" *)
  wire cbuf_p0_rd_sel_ram_b6c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:299" *)
  wire cbuf_p0_rd_sel_ram_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:96" *)
  wire cbuf_p0_rd_sel_ram_b7c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:300" *)
  wire cbuf_p0_rd_sel_ram_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:97" *)
  wire cbuf_p0_rd_sel_ram_b7c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:301" *)
  wire cbuf_p0_rd_sel_ram_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:98" *)
  wire cbuf_p0_rd_sel_ram_b8c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:302" *)
  wire cbuf_p0_rd_sel_ram_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:99" *)
  wire cbuf_p0_rd_sel_ram_b8c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:303" *)
  wire cbuf_p0_rd_sel_ram_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:100" *)
  wire cbuf_p0_rd_sel_ram_b9c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:304" *)
  wire cbuf_p0_rd_sel_ram_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:101" *)
  wire cbuf_p0_rd_sel_ram_b9c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:305" *)
  wire cbuf_p0_rd_sel_ram_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:306" *)
  reg cbuf_p0_rd_valid_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:102" *)
  wire [11:0] cbuf_p0_wr_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:307" *)
  reg [7:0] cbuf_p0_wr_addr_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:103" *)
  wire [3:0] cbuf_p0_wr_bank;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:104" *)
  wire cbuf_p0_wr_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:105" *)
  wire [511:0] cbuf_p0_wr_hi_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:308" *)
  reg [511:0] cbuf_p0_wr_hi_data_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:106" *)
  wire [511:0] cbuf_p0_wr_hi_data_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:107" *)
  wire cbuf_p0_wr_hi_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:108" *)
  wire cbuf_p0_wr_hi_en_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:109" *)
  wire [511:0] cbuf_p0_wr_lo_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:309" *)
  reg [511:0] cbuf_p0_wr_lo_data_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:110" *)
  wire [511:0] cbuf_p0_wr_lo_data_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:111" *)
  wire cbuf_p0_wr_lo_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:112" *)
  wire cbuf_p0_wr_lo_en_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:113" *)
  wire cbuf_p0_wr_sel_ram_b0c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:310" *)
  wire cbuf_p0_wr_sel_ram_b0c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:114" *)
  wire cbuf_p0_wr_sel_ram_b0c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:311" *)
  wire cbuf_p0_wr_sel_ram_b0c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:115" *)
  wire cbuf_p0_wr_sel_ram_b10c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:312" *)
  wire cbuf_p0_wr_sel_ram_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:116" *)
  wire cbuf_p0_wr_sel_ram_b10c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:313" *)
  wire cbuf_p0_wr_sel_ram_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:117" *)
  wire cbuf_p0_wr_sel_ram_b11c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:314" *)
  wire cbuf_p0_wr_sel_ram_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:118" *)
  wire cbuf_p0_wr_sel_ram_b11c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:315" *)
  wire cbuf_p0_wr_sel_ram_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:119" *)
  wire cbuf_p0_wr_sel_ram_b12c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:316" *)
  wire cbuf_p0_wr_sel_ram_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:120" *)
  wire cbuf_p0_wr_sel_ram_b12c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:317" *)
  wire cbuf_p0_wr_sel_ram_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:121" *)
  wire cbuf_p0_wr_sel_ram_b13c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:318" *)
  wire cbuf_p0_wr_sel_ram_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:122" *)
  wire cbuf_p0_wr_sel_ram_b13c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:319" *)
  wire cbuf_p0_wr_sel_ram_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:123" *)
  wire cbuf_p0_wr_sel_ram_b14c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:320" *)
  wire cbuf_p0_wr_sel_ram_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:124" *)
  wire cbuf_p0_wr_sel_ram_b14c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:321" *)
  wire cbuf_p0_wr_sel_ram_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:125" *)
  wire cbuf_p0_wr_sel_ram_b1c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:322" *)
  wire cbuf_p0_wr_sel_ram_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:126" *)
  wire cbuf_p0_wr_sel_ram_b1c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:323" *)
  wire cbuf_p0_wr_sel_ram_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:127" *)
  wire cbuf_p0_wr_sel_ram_b2c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:324" *)
  wire cbuf_p0_wr_sel_ram_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:128" *)
  wire cbuf_p0_wr_sel_ram_b2c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:325" *)
  wire cbuf_p0_wr_sel_ram_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:129" *)
  wire cbuf_p0_wr_sel_ram_b3c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:326" *)
  wire cbuf_p0_wr_sel_ram_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:130" *)
  wire cbuf_p0_wr_sel_ram_b3c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:327" *)
  wire cbuf_p0_wr_sel_ram_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:131" *)
  wire cbuf_p0_wr_sel_ram_b4c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:328" *)
  wire cbuf_p0_wr_sel_ram_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:132" *)
  wire cbuf_p0_wr_sel_ram_b4c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:329" *)
  wire cbuf_p0_wr_sel_ram_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:133" *)
  wire cbuf_p0_wr_sel_ram_b5c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:330" *)
  wire cbuf_p0_wr_sel_ram_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:134" *)
  wire cbuf_p0_wr_sel_ram_b5c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:331" *)
  wire cbuf_p0_wr_sel_ram_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:135" *)
  wire cbuf_p0_wr_sel_ram_b6c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:332" *)
  wire cbuf_p0_wr_sel_ram_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:136" *)
  wire cbuf_p0_wr_sel_ram_b6c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:333" *)
  wire cbuf_p0_wr_sel_ram_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:137" *)
  wire cbuf_p0_wr_sel_ram_b7c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:334" *)
  wire cbuf_p0_wr_sel_ram_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:138" *)
  wire cbuf_p0_wr_sel_ram_b7c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:335" *)
  wire cbuf_p0_wr_sel_ram_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:139" *)
  wire cbuf_p0_wr_sel_ram_b8c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:336" *)
  wire cbuf_p0_wr_sel_ram_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:140" *)
  wire cbuf_p0_wr_sel_ram_b8c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:337" *)
  wire cbuf_p0_wr_sel_ram_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:141" *)
  wire cbuf_p0_wr_sel_ram_b9c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:338" *)
  wire cbuf_p0_wr_sel_ram_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:142" *)
  wire cbuf_p0_wr_sel_ram_b9c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:339" *)
  wire cbuf_p0_wr_sel_ram_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:143" *)
  wire [11:0] cbuf_p1_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:144" *)
  wire [3:0] cbuf_p1_rd_bank;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:145" *)
  wire [511:0] cbuf_p1_rd_c0_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:340" *)
  reg [511:0] cbuf_p1_rd_c0_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:146" *)
  wire [511:0] cbuf_p1_rd_c0_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:341" *)
  wire cbuf_p1_rd_c0_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:147" *)
  wire cbuf_p1_rd_c0_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:148" *)
  wire [511:0] cbuf_p1_rd_c1_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:342" *)
  reg [511:0] cbuf_p1_rd_c1_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:149" *)
  wire [511:0] cbuf_p1_rd_c1_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:343" *)
  wire cbuf_p1_rd_c1_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:150" *)
  wire cbuf_p1_rd_c1_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:344" *)
  reg [1023:0] cbuf_p1_rd_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:345" *)
  wire [1023:0] cbuf_p1_rd_data_d4_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:346" *)
  reg [1023:0] cbuf_p1_rd_data_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:151" *)
  wire cbuf_p1_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:152" *)
  wire cbuf_p1_rd_en_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:153" *)
  wire cbuf_p1_rd_en_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:347" *)
  reg cbuf_p1_rd_en_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:154" *)
  wire cbuf_p1_rd_sel_ram_b10c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:348" *)
  wire cbuf_p1_rd_sel_ram_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:155" *)
  wire cbuf_p1_rd_sel_ram_b10c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:349" *)
  wire cbuf_p1_rd_sel_ram_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:156" *)
  wire cbuf_p1_rd_sel_ram_b11c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:350" *)
  wire cbuf_p1_rd_sel_ram_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:157" *)
  wire cbuf_p1_rd_sel_ram_b11c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:351" *)
  wire cbuf_p1_rd_sel_ram_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:158" *)
  wire cbuf_p1_rd_sel_ram_b12c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:352" *)
  wire cbuf_p1_rd_sel_ram_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:159" *)
  wire cbuf_p1_rd_sel_ram_b12c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:353" *)
  wire cbuf_p1_rd_sel_ram_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:160" *)
  wire cbuf_p1_rd_sel_ram_b13c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:354" *)
  wire cbuf_p1_rd_sel_ram_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:161" *)
  wire cbuf_p1_rd_sel_ram_b13c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:355" *)
  wire cbuf_p1_rd_sel_ram_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:162" *)
  wire cbuf_p1_rd_sel_ram_b14c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:356" *)
  wire cbuf_p1_rd_sel_ram_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:163" *)
  wire cbuf_p1_rd_sel_ram_b14c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:357" *)
  wire cbuf_p1_rd_sel_ram_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:164" *)
  wire cbuf_p1_rd_sel_ram_b15c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:358" *)
  wire cbuf_p1_rd_sel_ram_b15c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:165" *)
  wire cbuf_p1_rd_sel_ram_b15c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:359" *)
  wire cbuf_p1_rd_sel_ram_b15c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:166" *)
  wire cbuf_p1_rd_sel_ram_b1c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:360" *)
  wire cbuf_p1_rd_sel_ram_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:167" *)
  wire cbuf_p1_rd_sel_ram_b1c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:361" *)
  wire cbuf_p1_rd_sel_ram_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:168" *)
  wire cbuf_p1_rd_sel_ram_b2c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:362" *)
  wire cbuf_p1_rd_sel_ram_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:169" *)
  wire cbuf_p1_rd_sel_ram_b2c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:363" *)
  wire cbuf_p1_rd_sel_ram_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:170" *)
  wire cbuf_p1_rd_sel_ram_b3c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:364" *)
  wire cbuf_p1_rd_sel_ram_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:171" *)
  wire cbuf_p1_rd_sel_ram_b3c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:365" *)
  wire cbuf_p1_rd_sel_ram_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:172" *)
  wire cbuf_p1_rd_sel_ram_b4c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:366" *)
  wire cbuf_p1_rd_sel_ram_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:173" *)
  wire cbuf_p1_rd_sel_ram_b4c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:367" *)
  wire cbuf_p1_rd_sel_ram_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:174" *)
  wire cbuf_p1_rd_sel_ram_b5c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:368" *)
  wire cbuf_p1_rd_sel_ram_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:175" *)
  wire cbuf_p1_rd_sel_ram_b5c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:369" *)
  wire cbuf_p1_rd_sel_ram_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:176" *)
  wire cbuf_p1_rd_sel_ram_b6c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:370" *)
  wire cbuf_p1_rd_sel_ram_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:177" *)
  wire cbuf_p1_rd_sel_ram_b6c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:371" *)
  wire cbuf_p1_rd_sel_ram_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:178" *)
  wire cbuf_p1_rd_sel_ram_b7c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:372" *)
  wire cbuf_p1_rd_sel_ram_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:179" *)
  wire cbuf_p1_rd_sel_ram_b7c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:373" *)
  wire cbuf_p1_rd_sel_ram_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:180" *)
  wire cbuf_p1_rd_sel_ram_b8c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:374" *)
  wire cbuf_p1_rd_sel_ram_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:181" *)
  wire cbuf_p1_rd_sel_ram_b8c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:375" *)
  wire cbuf_p1_rd_sel_ram_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:182" *)
  wire cbuf_p1_rd_sel_ram_b9c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:376" *)
  wire cbuf_p1_rd_sel_ram_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:183" *)
  wire cbuf_p1_rd_sel_ram_b9c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:377" *)
  wire cbuf_p1_rd_sel_ram_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:378" *)
  reg cbuf_p1_rd_valid_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:184" *)
  wire [11:0] cbuf_p1_wr_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:379" *)
  reg [7:0] cbuf_p1_wr_addr_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:185" *)
  wire [3:0] cbuf_p1_wr_bank;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:186" *)
  wire [511:0] cbuf_p1_wr_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:187" *)
  wire cbuf_p1_wr_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:380" *)
  reg [511:0] cbuf_p1_wr_hi_data_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:188" *)
  wire [511:0] cbuf_p1_wr_hi_data_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:189" *)
  wire cbuf_p1_wr_hi_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:190" *)
  wire cbuf_p1_wr_hi_en_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:381" *)
  reg [511:0] cbuf_p1_wr_lo_data_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:191" *)
  wire [511:0] cbuf_p1_wr_lo_data_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:192" *)
  wire cbuf_p1_wr_lo_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:193" *)
  wire cbuf_p1_wr_lo_en_d1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:194" *)
  wire cbuf_p1_wr_sel_ram_b10c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:382" *)
  wire cbuf_p1_wr_sel_ram_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:195" *)
  wire cbuf_p1_wr_sel_ram_b10c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:383" *)
  wire cbuf_p1_wr_sel_ram_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:196" *)
  wire cbuf_p1_wr_sel_ram_b11c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:384" *)
  wire cbuf_p1_wr_sel_ram_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:197" *)
  wire cbuf_p1_wr_sel_ram_b11c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:385" *)
  wire cbuf_p1_wr_sel_ram_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:198" *)
  wire cbuf_p1_wr_sel_ram_b12c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:386" *)
  wire cbuf_p1_wr_sel_ram_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:199" *)
  wire cbuf_p1_wr_sel_ram_b12c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:387" *)
  wire cbuf_p1_wr_sel_ram_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:200" *)
  wire cbuf_p1_wr_sel_ram_b13c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:388" *)
  wire cbuf_p1_wr_sel_ram_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:201" *)
  wire cbuf_p1_wr_sel_ram_b13c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:389" *)
  wire cbuf_p1_wr_sel_ram_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:202" *)
  wire cbuf_p1_wr_sel_ram_b14c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:390" *)
  wire cbuf_p1_wr_sel_ram_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:203" *)
  wire cbuf_p1_wr_sel_ram_b14c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:391" *)
  wire cbuf_p1_wr_sel_ram_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:204" *)
  wire cbuf_p1_wr_sel_ram_b15c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:392" *)
  wire cbuf_p1_wr_sel_ram_b15c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:205" *)
  wire cbuf_p1_wr_sel_ram_b15c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:393" *)
  wire cbuf_p1_wr_sel_ram_b15c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:206" *)
  wire cbuf_p1_wr_sel_ram_b1c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:394" *)
  wire cbuf_p1_wr_sel_ram_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:207" *)
  wire cbuf_p1_wr_sel_ram_b1c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:395" *)
  wire cbuf_p1_wr_sel_ram_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:208" *)
  wire cbuf_p1_wr_sel_ram_b2c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:396" *)
  wire cbuf_p1_wr_sel_ram_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:209" *)
  wire cbuf_p1_wr_sel_ram_b2c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:397" *)
  wire cbuf_p1_wr_sel_ram_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:210" *)
  wire cbuf_p1_wr_sel_ram_b3c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:398" *)
  wire cbuf_p1_wr_sel_ram_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:211" *)
  wire cbuf_p1_wr_sel_ram_b3c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:399" *)
  wire cbuf_p1_wr_sel_ram_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:212" *)
  wire cbuf_p1_wr_sel_ram_b4c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:400" *)
  wire cbuf_p1_wr_sel_ram_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:213" *)
  wire cbuf_p1_wr_sel_ram_b4c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:401" *)
  wire cbuf_p1_wr_sel_ram_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:214" *)
  wire cbuf_p1_wr_sel_ram_b5c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:402" *)
  wire cbuf_p1_wr_sel_ram_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:215" *)
  wire cbuf_p1_wr_sel_ram_b5c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:403" *)
  wire cbuf_p1_wr_sel_ram_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:216" *)
  wire cbuf_p1_wr_sel_ram_b6c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:404" *)
  wire cbuf_p1_wr_sel_ram_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:217" *)
  wire cbuf_p1_wr_sel_ram_b6c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:405" *)
  wire cbuf_p1_wr_sel_ram_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:218" *)
  wire cbuf_p1_wr_sel_ram_b7c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:406" *)
  wire cbuf_p1_wr_sel_ram_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:219" *)
  wire cbuf_p1_wr_sel_ram_b7c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:407" *)
  wire cbuf_p1_wr_sel_ram_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:220" *)
  wire cbuf_p1_wr_sel_ram_b8c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:408" *)
  wire cbuf_p1_wr_sel_ram_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:221" *)
  wire cbuf_p1_wr_sel_ram_b8c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:409" *)
  wire cbuf_p1_wr_sel_ram_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:222" *)
  wire cbuf_p1_wr_sel_ram_b9c0_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:410" *)
  wire cbuf_p1_wr_sel_ram_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:223" *)
  wire cbuf_p1_wr_sel_ram_b9c1_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:411" *)
  wire cbuf_p1_wr_sel_ram_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:224" *)
  wire [7:0] cbuf_p2_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:225" *)
  wire [511:0] cbuf_p2_rd_c0_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:412" *)
  reg [511:0] cbuf_p2_rd_c0_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:226" *)
  wire [511:0] cbuf_p2_rd_c0_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:413" *)
  wire cbuf_p2_rd_c0_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:227" *)
  wire cbuf_p2_rd_c0_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:228" *)
  wire [511:0] cbuf_p2_rd_c1_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:414" *)
  reg [511:0] cbuf_p2_rd_c1_data_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:229" *)
  wire [511:0] cbuf_p2_rd_c1_data_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:415" *)
  wire cbuf_p2_rd_c1_valid_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:230" *)
  wire cbuf_p2_rd_c1_valid_d6_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:416" *)
  reg [1023:0] cbuf_p2_rd_data_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:417" *)
  wire [1023:0] cbuf_p2_rd_data_d4_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:418" *)
  reg [1023:0] cbuf_p2_rd_data_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:231" *)
  wire cbuf_p2_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:232" *)
  wire cbuf_p2_rd_en_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:233" *)
  wire cbuf_p2_rd_en_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:419" *)
  reg cbuf_p2_rd_en_d5;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:234" *)
  wire cbuf_p2_rd_sel_ram_b15c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:420" *)
  wire cbuf_p2_rd_sel_ram_b15c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:235" *)
  wire cbuf_p2_rd_sel_ram_b15c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:421" *)
  wire cbuf_p2_rd_sel_ram_b15c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:422" *)
  reg cbuf_p2_rd_valid_d6;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:423" *)
  reg [7:0] cbuf_ra_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:424" *)
  wire [7:0] cbuf_ra_b0c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:425" *)
  reg [7:0] cbuf_ra_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:426" *)
  wire [7:0] cbuf_ra_b0c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:427" *)
  reg [7:0] cbuf_ra_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:428" *)
  wire [7:0] cbuf_ra_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:429" *)
  reg [7:0] cbuf_ra_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:430" *)
  wire [7:0] cbuf_ra_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:431" *)
  reg [7:0] cbuf_ra_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:432" *)
  wire [7:0] cbuf_ra_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:433" *)
  reg [7:0] cbuf_ra_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:434" *)
  wire [7:0] cbuf_ra_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:435" *)
  reg [7:0] cbuf_ra_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:436" *)
  wire [7:0] cbuf_ra_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:437" *)
  reg [7:0] cbuf_ra_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:438" *)
  wire [7:0] cbuf_ra_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:439" *)
  reg [7:0] cbuf_ra_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:440" *)
  wire [7:0] cbuf_ra_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:441" *)
  reg [7:0] cbuf_ra_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:442" *)
  wire [7:0] cbuf_ra_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:443" *)
  reg [7:0] cbuf_ra_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:444" *)
  wire [7:0] cbuf_ra_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:445" *)
  reg [7:0] cbuf_ra_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:446" *)
  wire [7:0] cbuf_ra_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:447" *)
  reg [7:0] cbuf_ra_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:448" *)
  wire [7:0] cbuf_ra_b15c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:449" *)
  reg [7:0] cbuf_ra_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:450" *)
  wire [7:0] cbuf_ra_b15c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:451" *)
  reg [7:0] cbuf_ra_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:452" *)
  wire [7:0] cbuf_ra_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:453" *)
  reg [7:0] cbuf_ra_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:454" *)
  wire [7:0] cbuf_ra_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:455" *)
  reg [7:0] cbuf_ra_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:456" *)
  wire [7:0] cbuf_ra_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:457" *)
  reg [7:0] cbuf_ra_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:458" *)
  wire [7:0] cbuf_ra_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:459" *)
  reg [7:0] cbuf_ra_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:460" *)
  wire [7:0] cbuf_ra_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:461" *)
  reg [7:0] cbuf_ra_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:462" *)
  wire [7:0] cbuf_ra_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:463" *)
  reg [7:0] cbuf_ra_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:464" *)
  wire [7:0] cbuf_ra_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:465" *)
  reg [7:0] cbuf_ra_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:466" *)
  wire [7:0] cbuf_ra_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:467" *)
  reg [7:0] cbuf_ra_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:468" *)
  wire [7:0] cbuf_ra_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:469" *)
  reg [7:0] cbuf_ra_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:470" *)
  wire [7:0] cbuf_ra_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:471" *)
  reg [7:0] cbuf_ra_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:472" *)
  wire [7:0] cbuf_ra_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:473" *)
  reg [7:0] cbuf_ra_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:474" *)
  wire [7:0] cbuf_ra_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:475" *)
  reg [7:0] cbuf_ra_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:476" *)
  wire [7:0] cbuf_ra_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:477" *)
  reg [7:0] cbuf_ra_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:478" *)
  wire [7:0] cbuf_ra_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:479" *)
  reg [7:0] cbuf_ra_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:480" *)
  wire [7:0] cbuf_ra_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:481" *)
  reg [7:0] cbuf_ra_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:482" *)
  wire [7:0] cbuf_ra_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:483" *)
  reg [7:0] cbuf_ra_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:484" *)
  wire [7:0] cbuf_ra_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:485" *)
  reg [7:0] cbuf_ra_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:486" *)
  wire [7:0] cbuf_ra_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:487" *)
  reg [2:0] cbuf_rd_en_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:488" *)
  reg [2:0] cbuf_rd_en_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:489" *)
  reg [2:0] cbuf_rd_en_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:490" *)
  reg [2:0] cbuf_rd_en_d4;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:491" *)
  wire [61:0] cbuf_rd_sel_ram_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:492" *)
  wire [61:0] cbuf_rd_sel_ram_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:493" *)
  wire [61:0] cbuf_rd_sel_ram_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:236" *)
  wire [511:0] cbuf_rdat_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:494" *)
  reg [511:0] cbuf_rdat_b0c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:237" *)
  wire [511:0] cbuf_rdat_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:495" *)
  reg [511:0] cbuf_rdat_b0c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:238" *)
  wire [511:0] cbuf_rdat_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:496" *)
  reg [511:0] cbuf_rdat_b10c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:239" *)
  wire [511:0] cbuf_rdat_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:497" *)
  reg [511:0] cbuf_rdat_b10c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:240" *)
  wire [511:0] cbuf_rdat_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:498" *)
  reg [511:0] cbuf_rdat_b11c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:241" *)
  wire [511:0] cbuf_rdat_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:499" *)
  reg [511:0] cbuf_rdat_b11c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:242" *)
  wire [511:0] cbuf_rdat_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:500" *)
  reg [511:0] cbuf_rdat_b12c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:243" *)
  wire [511:0] cbuf_rdat_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:501" *)
  reg [511:0] cbuf_rdat_b12c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:244" *)
  wire [511:0] cbuf_rdat_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:502" *)
  reg [511:0] cbuf_rdat_b13c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:245" *)
  wire [511:0] cbuf_rdat_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:503" *)
  reg [511:0] cbuf_rdat_b13c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:246" *)
  wire [511:0] cbuf_rdat_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:504" *)
  reg [511:0] cbuf_rdat_b14c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:247" *)
  wire [511:0] cbuf_rdat_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:505" *)
  reg [511:0] cbuf_rdat_b14c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:248" *)
  wire [511:0] cbuf_rdat_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:506" *)
  reg [511:0] cbuf_rdat_b15c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:249" *)
  wire [511:0] cbuf_rdat_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:507" *)
  reg [511:0] cbuf_rdat_b15c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:250" *)
  wire [511:0] cbuf_rdat_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:508" *)
  reg [511:0] cbuf_rdat_b1c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:251" *)
  wire [511:0] cbuf_rdat_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:509" *)
  reg [511:0] cbuf_rdat_b1c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:252" *)
  wire [511:0] cbuf_rdat_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:510" *)
  reg [511:0] cbuf_rdat_b2c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:253" *)
  wire [511:0] cbuf_rdat_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:511" *)
  reg [511:0] cbuf_rdat_b2c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:254" *)
  wire [511:0] cbuf_rdat_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:512" *)
  reg [511:0] cbuf_rdat_b3c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:255" *)
  wire [511:0] cbuf_rdat_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:513" *)
  reg [511:0] cbuf_rdat_b3c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:256" *)
  wire [511:0] cbuf_rdat_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:514" *)
  reg [511:0] cbuf_rdat_b4c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:257" *)
  wire [511:0] cbuf_rdat_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:515" *)
  reg [511:0] cbuf_rdat_b4c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:258" *)
  wire [511:0] cbuf_rdat_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:516" *)
  reg [511:0] cbuf_rdat_b5c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:259" *)
  wire [511:0] cbuf_rdat_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:517" *)
  reg [511:0] cbuf_rdat_b5c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:260" *)
  wire [511:0] cbuf_rdat_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:518" *)
  reg [511:0] cbuf_rdat_b6c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:261" *)
  wire [511:0] cbuf_rdat_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:519" *)
  reg [511:0] cbuf_rdat_b6c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:262" *)
  wire [511:0] cbuf_rdat_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:520" *)
  reg [511:0] cbuf_rdat_b7c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:263" *)
  wire [511:0] cbuf_rdat_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:521" *)
  reg [511:0] cbuf_rdat_b7c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:264" *)
  wire [511:0] cbuf_rdat_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:522" *)
  reg [511:0] cbuf_rdat_b8c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:265" *)
  wire [511:0] cbuf_rdat_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:523" *)
  reg [511:0] cbuf_rdat_b8c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:266" *)
  wire [511:0] cbuf_rdat_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:524" *)
  reg [511:0] cbuf_rdat_b9c0_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:267" *)
  wire [511:0] cbuf_rdat_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:525" *)
  reg [511:0] cbuf_rdat_b9c1_d3;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:526" *)
  wire cbuf_re_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:527" *)
  wire cbuf_re_b0c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:528" *)
  wire cbuf_re_b0c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:529" *)
  reg cbuf_re_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:530" *)
  reg cbuf_re_b0c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:531" *)
  wire cbuf_re_b0c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:532" *)
  wire cbuf_re_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:533" *)
  wire cbuf_re_b10c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:534" *)
  wire cbuf_re_b10c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:535" *)
  reg cbuf_re_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:536" *)
  reg cbuf_re_b10c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:537" *)
  wire cbuf_re_b10c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:538" *)
  wire cbuf_re_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:539" *)
  wire cbuf_re_b11c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:540" *)
  wire cbuf_re_b11c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:541" *)
  reg cbuf_re_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:542" *)
  reg cbuf_re_b11c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:543" *)
  wire cbuf_re_b11c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:544" *)
  wire cbuf_re_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:545" *)
  wire cbuf_re_b12c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:546" *)
  wire cbuf_re_b12c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:547" *)
  reg cbuf_re_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:548" *)
  reg cbuf_re_b12c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:549" *)
  wire cbuf_re_b12c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:550" *)
  wire cbuf_re_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:551" *)
  wire cbuf_re_b13c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:552" *)
  wire cbuf_re_b13c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:553" *)
  reg cbuf_re_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:554" *)
  reg cbuf_re_b13c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:555" *)
  wire cbuf_re_b13c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:556" *)
  wire cbuf_re_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:557" *)
  wire cbuf_re_b14c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:558" *)
  wire cbuf_re_b14c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:559" *)
  reg cbuf_re_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:560" *)
  reg cbuf_re_b14c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:561" *)
  wire cbuf_re_b14c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:562" *)
  wire cbuf_re_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:563" *)
  wire cbuf_re_b15c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:564" *)
  wire cbuf_re_b15c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:565" *)
  reg cbuf_re_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:566" *)
  reg cbuf_re_b15c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:567" *)
  wire cbuf_re_b15c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:568" *)
  wire cbuf_re_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:569" *)
  wire cbuf_re_b1c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:570" *)
  wire cbuf_re_b1c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:571" *)
  reg cbuf_re_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:572" *)
  reg cbuf_re_b1c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:573" *)
  wire cbuf_re_b1c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:574" *)
  wire cbuf_re_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:575" *)
  wire cbuf_re_b2c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:576" *)
  wire cbuf_re_b2c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:577" *)
  reg cbuf_re_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:578" *)
  reg cbuf_re_b2c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:579" *)
  wire cbuf_re_b2c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:580" *)
  wire cbuf_re_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:581" *)
  wire cbuf_re_b3c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:582" *)
  wire cbuf_re_b3c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:583" *)
  reg cbuf_re_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:584" *)
  reg cbuf_re_b3c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:585" *)
  wire cbuf_re_b3c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:586" *)
  wire cbuf_re_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:587" *)
  wire cbuf_re_b4c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:588" *)
  wire cbuf_re_b4c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:589" *)
  reg cbuf_re_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:590" *)
  reg cbuf_re_b4c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:591" *)
  wire cbuf_re_b4c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:592" *)
  wire cbuf_re_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:593" *)
  wire cbuf_re_b5c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:594" *)
  wire cbuf_re_b5c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:595" *)
  reg cbuf_re_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:596" *)
  reg cbuf_re_b5c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:597" *)
  wire cbuf_re_b5c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:598" *)
  wire cbuf_re_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:599" *)
  wire cbuf_re_b6c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:600" *)
  wire cbuf_re_b6c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:601" *)
  reg cbuf_re_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:602" *)
  reg cbuf_re_b6c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:603" *)
  wire cbuf_re_b6c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:604" *)
  wire cbuf_re_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:605" *)
  wire cbuf_re_b7c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:606" *)
  wire cbuf_re_b7c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:607" *)
  reg cbuf_re_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:608" *)
  reg cbuf_re_b7c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:609" *)
  wire cbuf_re_b7c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:610" *)
  wire cbuf_re_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:611" *)
  wire cbuf_re_b8c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:612" *)
  wire cbuf_re_b8c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:613" *)
  reg cbuf_re_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:614" *)
  reg cbuf_re_b8c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:615" *)
  wire cbuf_re_b8c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:616" *)
  wire cbuf_re_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:617" *)
  wire cbuf_re_b9c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:618" *)
  wire cbuf_re_b9c0_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:619" *)
  reg cbuf_re_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:620" *)
  reg cbuf_re_b9c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:621" *)
  wire cbuf_re_b9c1_w;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:622" *)
  wire [7:0] cbuf_wa_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:623" *)
  reg [7:0] cbuf_wa_b0c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:624" *)
  wire [7:0] cbuf_wa_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:625" *)
  reg [7:0] cbuf_wa_b0c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:626" *)
  wire [7:0] cbuf_wa_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:627" *)
  reg [7:0] cbuf_wa_b10c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:628" *)
  wire [7:0] cbuf_wa_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:629" *)
  reg [7:0] cbuf_wa_b10c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:630" *)
  wire [7:0] cbuf_wa_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:631" *)
  reg [7:0] cbuf_wa_b11c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:632" *)
  wire [7:0] cbuf_wa_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:633" *)
  reg [7:0] cbuf_wa_b11c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:634" *)
  wire [7:0] cbuf_wa_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:635" *)
  reg [7:0] cbuf_wa_b12c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:636" *)
  wire [7:0] cbuf_wa_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:637" *)
  reg [7:0] cbuf_wa_b12c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:638" *)
  wire [7:0] cbuf_wa_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:639" *)
  reg [7:0] cbuf_wa_b13c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:640" *)
  wire [7:0] cbuf_wa_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:641" *)
  reg [7:0] cbuf_wa_b13c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:642" *)
  wire [7:0] cbuf_wa_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:643" *)
  reg [7:0] cbuf_wa_b14c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:644" *)
  wire [7:0] cbuf_wa_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:645" *)
  reg [7:0] cbuf_wa_b14c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:646" *)
  wire [7:0] cbuf_wa_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:647" *)
  reg [7:0] cbuf_wa_b15c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:648" *)
  wire [7:0] cbuf_wa_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:649" *)
  reg [7:0] cbuf_wa_b15c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:650" *)
  wire [7:0] cbuf_wa_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:651" *)
  reg [7:0] cbuf_wa_b1c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:652" *)
  wire [7:0] cbuf_wa_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:653" *)
  reg [7:0] cbuf_wa_b1c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:654" *)
  wire [7:0] cbuf_wa_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:655" *)
  reg [7:0] cbuf_wa_b2c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:656" *)
  wire [7:0] cbuf_wa_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:657" *)
  reg [7:0] cbuf_wa_b2c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:658" *)
  wire [7:0] cbuf_wa_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:659" *)
  reg [7:0] cbuf_wa_b3c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:660" *)
  wire [7:0] cbuf_wa_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:661" *)
  reg [7:0] cbuf_wa_b3c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:662" *)
  wire [7:0] cbuf_wa_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:663" *)
  reg [7:0] cbuf_wa_b4c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:664" *)
  wire [7:0] cbuf_wa_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:665" *)
  reg [7:0] cbuf_wa_b4c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:666" *)
  wire [7:0] cbuf_wa_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:667" *)
  reg [7:0] cbuf_wa_b5c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:668" *)
  wire [7:0] cbuf_wa_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:669" *)
  reg [7:0] cbuf_wa_b5c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:670" *)
  wire [7:0] cbuf_wa_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:671" *)
  reg [7:0] cbuf_wa_b6c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:672" *)
  wire [7:0] cbuf_wa_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:673" *)
  reg [7:0] cbuf_wa_b6c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:674" *)
  wire [7:0] cbuf_wa_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:675" *)
  reg [7:0] cbuf_wa_b7c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:676" *)
  wire [7:0] cbuf_wa_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:677" *)
  reg [7:0] cbuf_wa_b7c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:678" *)
  wire [7:0] cbuf_wa_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:679" *)
  reg [7:0] cbuf_wa_b8c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:680" *)
  wire [7:0] cbuf_wa_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:681" *)
  reg [7:0] cbuf_wa_b8c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:682" *)
  wire [7:0] cbuf_wa_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:683" *)
  reg [7:0] cbuf_wa_b9c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:684" *)
  wire [7:0] cbuf_wa_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:685" *)
  reg [7:0] cbuf_wa_b9c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:686" *)
  wire [511:0] cbuf_wdat_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:687" *)
  reg [511:0] cbuf_wdat_b0c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:688" *)
  wire [511:0] cbuf_wdat_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:689" *)
  reg [511:0] cbuf_wdat_b0c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:690" *)
  wire [511:0] cbuf_wdat_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:691" *)
  reg [511:0] cbuf_wdat_b10c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:692" *)
  wire [511:0] cbuf_wdat_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:693" *)
  reg [511:0] cbuf_wdat_b10c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:694" *)
  wire [511:0] cbuf_wdat_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:695" *)
  reg [511:0] cbuf_wdat_b11c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:696" *)
  wire [511:0] cbuf_wdat_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:697" *)
  reg [511:0] cbuf_wdat_b11c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:698" *)
  wire [511:0] cbuf_wdat_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:699" *)
  reg [511:0] cbuf_wdat_b12c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:700" *)
  wire [511:0] cbuf_wdat_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:701" *)
  reg [511:0] cbuf_wdat_b12c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:702" *)
  wire [511:0] cbuf_wdat_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:703" *)
  reg [511:0] cbuf_wdat_b13c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:704" *)
  wire [511:0] cbuf_wdat_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:705" *)
  reg [511:0] cbuf_wdat_b13c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:706" *)
  wire [511:0] cbuf_wdat_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:707" *)
  reg [511:0] cbuf_wdat_b14c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:708" *)
  wire [511:0] cbuf_wdat_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:709" *)
  reg [511:0] cbuf_wdat_b14c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:710" *)
  wire [511:0] cbuf_wdat_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:711" *)
  reg [511:0] cbuf_wdat_b15c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:712" *)
  wire [511:0] cbuf_wdat_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:713" *)
  reg [511:0] cbuf_wdat_b15c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:714" *)
  wire [511:0] cbuf_wdat_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:715" *)
  reg [511:0] cbuf_wdat_b1c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:716" *)
  wire [511:0] cbuf_wdat_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:717" *)
  reg [511:0] cbuf_wdat_b1c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:718" *)
  wire [511:0] cbuf_wdat_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:719" *)
  reg [511:0] cbuf_wdat_b2c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:720" *)
  wire [511:0] cbuf_wdat_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:721" *)
  reg [511:0] cbuf_wdat_b2c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:722" *)
  wire [511:0] cbuf_wdat_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:723" *)
  reg [511:0] cbuf_wdat_b3c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:724" *)
  wire [511:0] cbuf_wdat_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:725" *)
  reg [511:0] cbuf_wdat_b3c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:726" *)
  wire [511:0] cbuf_wdat_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:727" *)
  reg [511:0] cbuf_wdat_b4c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:728" *)
  wire [511:0] cbuf_wdat_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:729" *)
  reg [511:0] cbuf_wdat_b4c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:730" *)
  wire [511:0] cbuf_wdat_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:731" *)
  reg [511:0] cbuf_wdat_b5c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:732" *)
  wire [511:0] cbuf_wdat_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:733" *)
  reg [511:0] cbuf_wdat_b5c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:734" *)
  wire [511:0] cbuf_wdat_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:735" *)
  reg [511:0] cbuf_wdat_b6c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:736" *)
  wire [511:0] cbuf_wdat_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:737" *)
  reg [511:0] cbuf_wdat_b6c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:738" *)
  wire [511:0] cbuf_wdat_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:739" *)
  reg [511:0] cbuf_wdat_b7c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:740" *)
  wire [511:0] cbuf_wdat_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:741" *)
  reg [511:0] cbuf_wdat_b7c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:742" *)
  wire [511:0] cbuf_wdat_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:743" *)
  reg [511:0] cbuf_wdat_b8c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:744" *)
  wire [511:0] cbuf_wdat_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:745" *)
  reg [511:0] cbuf_wdat_b8c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:746" *)
  wire [511:0] cbuf_wdat_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:747" *)
  reg [511:0] cbuf_wdat_b9c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:748" *)
  wire [511:0] cbuf_wdat_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:749" *)
  reg [511:0] cbuf_wdat_b9c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:750" *)
  reg cbuf_we_b0c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:751" *)
  reg cbuf_we_b0c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:752" *)
  reg cbuf_we_b0c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:753" *)
  reg cbuf_we_b0c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:754" *)
  reg cbuf_we_b10c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:755" *)
  reg cbuf_we_b10c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:756" *)
  reg cbuf_we_b10c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:757" *)
  reg cbuf_we_b10c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:758" *)
  reg cbuf_we_b11c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:759" *)
  reg cbuf_we_b11c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:760" *)
  reg cbuf_we_b11c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:761" *)
  reg cbuf_we_b11c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:762" *)
  reg cbuf_we_b12c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:763" *)
  reg cbuf_we_b12c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:764" *)
  reg cbuf_we_b12c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:765" *)
  reg cbuf_we_b12c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:766" *)
  reg cbuf_we_b13c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:767" *)
  reg cbuf_we_b13c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:768" *)
  reg cbuf_we_b13c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:769" *)
  reg cbuf_we_b13c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:770" *)
  reg cbuf_we_b14c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:771" *)
  reg cbuf_we_b14c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:772" *)
  reg cbuf_we_b14c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:773" *)
  reg cbuf_we_b14c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:774" *)
  reg cbuf_we_b15c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:775" *)
  reg cbuf_we_b15c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:776" *)
  reg cbuf_we_b15c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:777" *)
  reg cbuf_we_b15c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:778" *)
  reg cbuf_we_b1c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:779" *)
  reg cbuf_we_b1c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:780" *)
  reg cbuf_we_b1c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:781" *)
  reg cbuf_we_b1c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:782" *)
  reg cbuf_we_b2c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:783" *)
  reg cbuf_we_b2c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:784" *)
  reg cbuf_we_b2c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:785" *)
  reg cbuf_we_b2c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:786" *)
  reg cbuf_we_b3c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:787" *)
  reg cbuf_we_b3c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:788" *)
  reg cbuf_we_b3c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:789" *)
  reg cbuf_we_b3c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:790" *)
  reg cbuf_we_b4c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:791" *)
  reg cbuf_we_b4c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:792" *)
  reg cbuf_we_b4c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:793" *)
  reg cbuf_we_b4c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:794" *)
  reg cbuf_we_b5c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:795" *)
  reg cbuf_we_b5c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:796" *)
  reg cbuf_we_b5c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:797" *)
  reg cbuf_we_b5c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:798" *)
  reg cbuf_we_b6c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:799" *)
  reg cbuf_we_b6c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:800" *)
  reg cbuf_we_b6c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:801" *)
  reg cbuf_we_b6c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:802" *)
  reg cbuf_we_b7c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:803" *)
  reg cbuf_we_b7c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:804" *)
  reg cbuf_we_b7c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:805" *)
  reg cbuf_we_b7c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:806" *)
  reg cbuf_we_b8c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:807" *)
  reg cbuf_we_b8c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:808" *)
  reg cbuf_we_b8c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:809" *)
  reg cbuf_we_b8c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:810" *)
  reg cbuf_we_b9c0;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:811" *)
  reg cbuf_we_b9c0_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:812" *)
  reg cbuf_we_b9c1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:813" *)
  reg cbuf_we_b9c1_d2;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:814" *)
  reg [59:0] cbuf_wr_sel_ram_d1;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:42" *)
  input [11:0] cdma2buf_dat_wr_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:44" *)
  input [1023:0] cdma2buf_dat_wr_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:41" *)
  input cdma2buf_dat_wr_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:43" *)
  input [1:0] cdma2buf_dat_wr_hsel;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:46" *)
  input [11:0] cdma2buf_wt_wr_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:48" *)
  input [511:0] cdma2buf_wt_wr_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:45" *)
  input cdma2buf_wt_wr_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:47" *)
  input cdma2buf_wt_wr_hsel;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:38" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:39" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:40" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:50" *)
  input [11:0] sc2buf_dat_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:52" *)
  output [1023:0] sc2buf_dat_rd_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:49" *)
  input sc2buf_dat_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:51" *)
  output sc2buf_dat_rd_valid;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:58" *)
  input [7:0] sc2buf_wmb_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:60" *)
  output [1023:0] sc2buf_wmb_rd_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:57" *)
  input sc2buf_wmb_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:59" *)
  output sc2buf_wmb_rd_valid;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:54" *)
  input [11:0] sc2buf_wt_rd_addr;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:56" *)
  output [1023:0] sc2buf_wt_rd_data;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:53" *)
  input sc2buf_wt_rd_en;
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:55" *)
  output sc2buf_wt_rd_valid;
  assign cbuf_wa_b0c0 = { cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1693" *) cbuf_p0_wr_addr_d1;
  assign cbuf_wdat_b0c0 = { cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59], cbuf_wr_sel_ram_d1[59] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1694" *) cbuf_p0_wr_lo_data_d1;
  assign cbuf_wa_b0c1 = { cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1701" *) cbuf_p0_wr_addr_d1;
  assign cbuf_wdat_b0c1 = { cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58], cbuf_wr_sel_ram_d1[58] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1702" *) cbuf_p0_wr_hi_data_d1;
  assign _0180_ = { cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1712" *) cbuf_p0_wr_addr_d1;
  assign _0181_ = { cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1713" *) cbuf_p1_wr_addr_d1;
  assign _0182_ = { cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57], cbuf_wr_sel_ram_d1[57] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1714" *) cbuf_p0_wr_lo_data_d1;
  assign _0183_ = { cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29], cbuf_wr_sel_ram_d1[29] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1715" *) cbuf_p1_wr_lo_data_d1;
  assign _0184_ = { cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1725" *) cbuf_p0_wr_addr_d1;
  assign _0185_ = { cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1726" *) cbuf_p1_wr_addr_d1;
  assign _0186_ = { cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56], cbuf_wr_sel_ram_d1[56] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1727" *) cbuf_p0_wr_hi_data_d1;
  assign _0187_ = { cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28], cbuf_wr_sel_ram_d1[28] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1728" *) cbuf_p1_wr_hi_data_d1;
  assign _0188_ = { cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1738" *) cbuf_p0_wr_addr_d1;
  assign _0189_ = { cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1739" *) cbuf_p1_wr_addr_d1;
  assign _0190_ = { cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55], cbuf_wr_sel_ram_d1[55] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1740" *) cbuf_p0_wr_lo_data_d1;
  assign _0191_ = { cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27], cbuf_wr_sel_ram_d1[27] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1741" *) cbuf_p1_wr_lo_data_d1;
  assign _0192_ = { cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1751" *) cbuf_p0_wr_addr_d1;
  assign _0193_ = { cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1752" *) cbuf_p1_wr_addr_d1;
  assign _0194_ = { cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54], cbuf_wr_sel_ram_d1[54] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1753" *) cbuf_p0_wr_hi_data_d1;
  assign _0195_ = { cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26], cbuf_wr_sel_ram_d1[26] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1754" *) cbuf_p1_wr_hi_data_d1;
  assign _0196_ = { cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1764" *) cbuf_p0_wr_addr_d1;
  assign _0197_ = { cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1765" *) cbuf_p1_wr_addr_d1;
  assign _0198_ = { cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53], cbuf_wr_sel_ram_d1[53] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1766" *) cbuf_p0_wr_lo_data_d1;
  assign _0199_ = { cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25], cbuf_wr_sel_ram_d1[25] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1767" *) cbuf_p1_wr_lo_data_d1;
  assign _0200_ = { cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1777" *) cbuf_p0_wr_addr_d1;
  assign _0201_ = { cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1778" *) cbuf_p1_wr_addr_d1;
  assign _0202_ = { cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52], cbuf_wr_sel_ram_d1[52] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1779" *) cbuf_p0_wr_hi_data_d1;
  assign _0203_ = { cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24], cbuf_wr_sel_ram_d1[24] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1780" *) cbuf_p1_wr_hi_data_d1;
  assign _0204_ = { cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1790" *) cbuf_p0_wr_addr_d1;
  assign _0205_ = { cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1791" *) cbuf_p1_wr_addr_d1;
  assign _0206_ = { cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51], cbuf_wr_sel_ram_d1[51] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1792" *) cbuf_p0_wr_lo_data_d1;
  assign _0207_ = { cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23], cbuf_wr_sel_ram_d1[23] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1793" *) cbuf_p1_wr_lo_data_d1;
  assign _0208_ = { cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1803" *) cbuf_p0_wr_addr_d1;
  assign _0209_ = { cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1804" *) cbuf_p1_wr_addr_d1;
  assign _0210_ = { cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50], cbuf_wr_sel_ram_d1[50] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1805" *) cbuf_p0_wr_hi_data_d1;
  assign _0211_ = { cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22], cbuf_wr_sel_ram_d1[22] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1806" *) cbuf_p1_wr_hi_data_d1;
  assign _0212_ = { cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1816" *) cbuf_p0_wr_addr_d1;
  assign _0213_ = { cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1817" *) cbuf_p1_wr_addr_d1;
  assign _0214_ = { cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49], cbuf_wr_sel_ram_d1[49] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1818" *) cbuf_p0_wr_lo_data_d1;
  assign _0215_ = { cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21], cbuf_wr_sel_ram_d1[21] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1819" *) cbuf_p1_wr_lo_data_d1;
  assign _0216_ = { cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1829" *) cbuf_p0_wr_addr_d1;
  assign _0217_ = { cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1830" *) cbuf_p1_wr_addr_d1;
  assign _0218_ = { cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48], cbuf_wr_sel_ram_d1[48] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1831" *) cbuf_p0_wr_hi_data_d1;
  assign _0219_ = { cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20], cbuf_wr_sel_ram_d1[20] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1832" *) cbuf_p1_wr_hi_data_d1;
  assign _0220_ = { cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1842" *) cbuf_p0_wr_addr_d1;
  assign _0221_ = { cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1843" *) cbuf_p1_wr_addr_d1;
  assign _0222_ = { cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47], cbuf_wr_sel_ram_d1[47] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1844" *) cbuf_p0_wr_lo_data_d1;
  assign _0223_ = { cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19], cbuf_wr_sel_ram_d1[19] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1845" *) cbuf_p1_wr_lo_data_d1;
  assign _0224_ = { cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1855" *) cbuf_p0_wr_addr_d1;
  assign _0225_ = { cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1856" *) cbuf_p1_wr_addr_d1;
  assign _0226_ = { cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46], cbuf_wr_sel_ram_d1[46] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1857" *) cbuf_p0_wr_hi_data_d1;
  assign _0227_ = { cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18], cbuf_wr_sel_ram_d1[18] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1858" *) cbuf_p1_wr_hi_data_d1;
  assign _0228_ = { cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1868" *) cbuf_p0_wr_addr_d1;
  assign _0229_ = { cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1869" *) cbuf_p1_wr_addr_d1;
  assign _0230_ = { cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45], cbuf_wr_sel_ram_d1[45] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1870" *) cbuf_p0_wr_lo_data_d1;
  assign _0231_ = { cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17], cbuf_wr_sel_ram_d1[17] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1871" *) cbuf_p1_wr_lo_data_d1;
  assign _0232_ = { cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1881" *) cbuf_p0_wr_addr_d1;
  assign _0233_ = { cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1882" *) cbuf_p1_wr_addr_d1;
  assign _0234_ = { cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44], cbuf_wr_sel_ram_d1[44] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1883" *) cbuf_p0_wr_hi_data_d1;
  assign _0235_ = { cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16], cbuf_wr_sel_ram_d1[16] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1884" *) cbuf_p1_wr_hi_data_d1;
  assign _0236_ = { cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1894" *) cbuf_p0_wr_addr_d1;
  assign _0237_ = { cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1895" *) cbuf_p1_wr_addr_d1;
  assign _0238_ = { cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43], cbuf_wr_sel_ram_d1[43] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1896" *) cbuf_p0_wr_lo_data_d1;
  assign _0239_ = { cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15], cbuf_wr_sel_ram_d1[15] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1897" *) cbuf_p1_wr_lo_data_d1;
  assign _0240_ = { cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1907" *) cbuf_p0_wr_addr_d1;
  assign _0241_ = { cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1908" *) cbuf_p1_wr_addr_d1;
  assign _0242_ = { cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42], cbuf_wr_sel_ram_d1[42] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1909" *) cbuf_p0_wr_hi_data_d1;
  assign _0243_ = { cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14], cbuf_wr_sel_ram_d1[14] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1910" *) cbuf_p1_wr_hi_data_d1;
  assign _0244_ = { cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1920" *) cbuf_p0_wr_addr_d1;
  assign _0245_ = { cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1921" *) cbuf_p1_wr_addr_d1;
  assign _0246_ = { cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41], cbuf_wr_sel_ram_d1[41] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1922" *) cbuf_p0_wr_lo_data_d1;
  assign _0247_ = { cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13], cbuf_wr_sel_ram_d1[13] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1923" *) cbuf_p1_wr_lo_data_d1;
  assign _0248_ = { cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1933" *) cbuf_p0_wr_addr_d1;
  assign _0249_ = { cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1934" *) cbuf_p1_wr_addr_d1;
  assign _0250_ = { cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40], cbuf_wr_sel_ram_d1[40] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1935" *) cbuf_p0_wr_hi_data_d1;
  assign _0251_ = { cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12], cbuf_wr_sel_ram_d1[12] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1936" *) cbuf_p1_wr_hi_data_d1;
  assign _0252_ = { cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1946" *) cbuf_p0_wr_addr_d1;
  assign _0253_ = { cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1947" *) cbuf_p1_wr_addr_d1;
  assign _0254_ = { cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39], cbuf_wr_sel_ram_d1[39] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1948" *) cbuf_p0_wr_lo_data_d1;
  assign _0255_ = { cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11], cbuf_wr_sel_ram_d1[11] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1949" *) cbuf_p1_wr_lo_data_d1;
  assign _0256_ = { cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1959" *) cbuf_p0_wr_addr_d1;
  assign _0257_ = { cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1960" *) cbuf_p1_wr_addr_d1;
  assign _0258_ = { cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38], cbuf_wr_sel_ram_d1[38] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1961" *) cbuf_p0_wr_hi_data_d1;
  assign _0259_ = { cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10], cbuf_wr_sel_ram_d1[10] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1962" *) cbuf_p1_wr_hi_data_d1;
  assign _0260_ = { cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1972" *) cbuf_p0_wr_addr_d1;
  assign _0261_ = { cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1973" *) cbuf_p1_wr_addr_d1;
  assign _0262_ = { cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37], cbuf_wr_sel_ram_d1[37] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1974" *) cbuf_p0_wr_lo_data_d1;
  assign _0263_ = { cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9], cbuf_wr_sel_ram_d1[9] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1975" *) cbuf_p1_wr_lo_data_d1;
  assign _0264_ = { cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1985" *) cbuf_p0_wr_addr_d1;
  assign _0265_ = { cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1986" *) cbuf_p1_wr_addr_d1;
  assign _0266_ = { cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36], cbuf_wr_sel_ram_d1[36] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1987" *) cbuf_p0_wr_hi_data_d1;
  assign _0267_ = { cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8], cbuf_wr_sel_ram_d1[8] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1988" *) cbuf_p1_wr_hi_data_d1;
  assign _0268_ = { cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1998" *) cbuf_p0_wr_addr_d1;
  assign _0269_ = { cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1999" *) cbuf_p1_wr_addr_d1;
  assign _0270_ = { cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35], cbuf_wr_sel_ram_d1[35] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2000" *) cbuf_p0_wr_lo_data_d1;
  assign _0271_ = { cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7], cbuf_wr_sel_ram_d1[7] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2001" *) cbuf_p1_wr_lo_data_d1;
  assign _0272_ = { cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2011" *) cbuf_p0_wr_addr_d1;
  assign _0273_ = { cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2012" *) cbuf_p1_wr_addr_d1;
  assign _0274_ = { cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34], cbuf_wr_sel_ram_d1[34] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2013" *) cbuf_p0_wr_hi_data_d1;
  assign _0275_ = { cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6], cbuf_wr_sel_ram_d1[6] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2014" *) cbuf_p1_wr_hi_data_d1;
  assign _0276_ = { cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2024" *) cbuf_p0_wr_addr_d1;
  assign _0277_ = { cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2025" *) cbuf_p1_wr_addr_d1;
  assign _0278_ = { cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33], cbuf_wr_sel_ram_d1[33] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2026" *) cbuf_p0_wr_lo_data_d1;
  assign _0279_ = { cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5], cbuf_wr_sel_ram_d1[5] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2027" *) cbuf_p1_wr_lo_data_d1;
  assign _0280_ = { cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2037" *) cbuf_p0_wr_addr_d1;
  assign _0281_ = { cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2038" *) cbuf_p1_wr_addr_d1;
  assign _0282_ = { cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32], cbuf_wr_sel_ram_d1[32] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2039" *) cbuf_p0_wr_hi_data_d1;
  assign _0283_ = { cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4], cbuf_wr_sel_ram_d1[4] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2040" *) cbuf_p1_wr_hi_data_d1;
  assign _0284_ = { cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2050" *) cbuf_p0_wr_addr_d1;
  assign _0285_ = { cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2051" *) cbuf_p1_wr_addr_d1;
  assign _0286_ = { cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31], cbuf_wr_sel_ram_d1[31] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2052" *) cbuf_p0_wr_lo_data_d1;
  assign _0287_ = { cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3], cbuf_wr_sel_ram_d1[3] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2053" *) cbuf_p1_wr_lo_data_d1;
  assign _0288_ = { cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2063" *) cbuf_p0_wr_addr_d1;
  assign _0289_ = { cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2064" *) cbuf_p1_wr_addr_d1;
  assign _0290_ = { cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30], cbuf_wr_sel_ram_d1[30] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2065" *) cbuf_p0_wr_hi_data_d1;
  assign _0291_ = { cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2], cbuf_wr_sel_ram_d1[2] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2066" *) cbuf_p1_wr_hi_data_d1;
  assign cbuf_wa_b15c0 = { cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2073" *) cbuf_p1_wr_addr_d1;
  assign cbuf_wdat_b15c0 = { cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1], cbuf_wr_sel_ram_d1[1] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2074" *) cbuf_p1_wr_lo_data_d1;
  assign cbuf_wa_b15c1 = { cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2081" *) cbuf_p1_wr_addr_d1;
  assign cbuf_wdat_b15c1 = { cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0], cbuf_wr_sel_ram_d1[0] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2082" *) cbuf_p1_wr_hi_data_d1;
  assign cbuf_ra_b0c0_w = { cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b0c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3912" *) sc2buf_dat_rd_addr[7:0];
  assign _0292_ = { cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3926" *) sc2buf_dat_rd_addr[7:0];
  assign _0293_ = { cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3927" *) sc2buf_wt_rd_addr[7:0];
  assign _0294_ = { cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3953" *) sc2buf_dat_rd_addr[7:0];
  assign _0295_ = { cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3954" *) sc2buf_wt_rd_addr[7:0];
  assign _0296_ = { cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3962" *) sc2buf_dat_rd_addr[7:0];
  assign _0297_ = { cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3963" *) sc2buf_wt_rd_addr[7:0];
  assign _0298_ = { cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3980" *) sc2buf_dat_rd_addr[7:0];
  assign _0299_ = { cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3981" *) sc2buf_wt_rd_addr[7:0];
  assign _0300_ = { cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3998" *) sc2buf_dat_rd_addr[7:0];
  assign _0301_ = { cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3999" *) sc2buf_wt_rd_addr[7:0];
  assign _0302_ = { cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4016" *) sc2buf_dat_rd_addr[7:0];
  assign _0303_ = { cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4017" *) sc2buf_wt_rd_addr[7:0];
  assign _0304_ = { cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4034" *) sc2buf_dat_rd_addr[7:0];
  assign _0305_ = { cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4035" *) sc2buf_wt_rd_addr[7:0];
  assign _0306_ = { cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4052" *) sc2buf_dat_rd_addr[7:0];
  assign _0307_ = { cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4053" *) sc2buf_wt_rd_addr[7:0];
  assign _0308_ = { cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4070" *) sc2buf_dat_rd_addr[7:0];
  assign _0309_ = { cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4071" *) sc2buf_wt_rd_addr[7:0];
  assign _0310_ = { cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4088" *) sc2buf_dat_rd_addr[7:0];
  assign _0311_ = { cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4089" *) sc2buf_wt_rd_addr[7:0];
  assign _0312_ = { cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4106" *) sc2buf_dat_rd_addr[7:0];
  assign _0313_ = { cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4107" *) sc2buf_wt_rd_addr[7:0];
  assign _0314_ = { cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4124" *) sc2buf_dat_rd_addr[7:0];
  assign _0315_ = { cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4125" *) sc2buf_wt_rd_addr[7:0];
  assign _0316_ = { cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4142" *) sc2buf_dat_rd_addr[7:0];
  assign _0317_ = { cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4143" *) sc2buf_wt_rd_addr[7:0];
  assign _0318_ = { cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4160" *) sc2buf_dat_rd_addr[7:0];
  assign _0319_ = { cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4161" *) sc2buf_wt_rd_addr[7:0];
  assign _0320_ = { cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4178" *) sc2buf_wt_rd_addr[7:0];
  assign _0321_ = { sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4179" *) sc2buf_wmb_rd_addr;
  assign _0322_ = { cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60], cbuf_rd_sel_ram_d3[60] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5525" *) { cbuf_rdat_b0c0_d3, cbuf_rdat_b0c1_d3 };
  assign _0323_ = { cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59], cbuf_rd_sel_ram_d3[59:58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58], cbuf_rd_sel_ram_d3[58] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5526" *) { cbuf_rdat_b1c0_d3, cbuf_rdat_b1c1_d3 };
  assign _0324_ = { cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57], cbuf_rd_sel_ram_d3[57:56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56], cbuf_rd_sel_ram_d3[56] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5527" *) { cbuf_rdat_b2c0_d3, cbuf_rdat_b2c1_d3 };
  assign _0325_ = { cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55], cbuf_rd_sel_ram_d3[55:54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54], cbuf_rd_sel_ram_d3[54] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5528" *) { cbuf_rdat_b3c0_d3, cbuf_rdat_b3c1_d3 };
  assign _0326_ = { cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53], cbuf_rd_sel_ram_d3[53:52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52], cbuf_rd_sel_ram_d3[52] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5529" *) { cbuf_rdat_b4c0_d3, cbuf_rdat_b4c1_d3 };
  assign _0327_ = { cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51], cbuf_rd_sel_ram_d3[51:50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50], cbuf_rd_sel_ram_d3[50] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5530" *) { cbuf_rdat_b5c0_d3, cbuf_rdat_b5c1_d3 };
  assign _0328_ = { cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49], cbuf_rd_sel_ram_d3[49:48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48], cbuf_rd_sel_ram_d3[48] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5531" *) { cbuf_rdat_b6c0_d3, cbuf_rdat_b6c1_d3 };
  assign _0329_ = { cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47], cbuf_rd_sel_ram_d3[47:46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46], cbuf_rd_sel_ram_d3[46] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5532" *) { cbuf_rdat_b7c0_d3, cbuf_rdat_b7c1_d3 };
  assign _0330_ = { cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45], cbuf_rd_sel_ram_d3[45:44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44], cbuf_rd_sel_ram_d3[44] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5533" *) { cbuf_rdat_b8c0_d3, cbuf_rdat_b8c1_d3 };
  assign _0331_ = { cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43], cbuf_rd_sel_ram_d3[43:42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42], cbuf_rd_sel_ram_d3[42] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5534" *) { cbuf_rdat_b9c0_d3, cbuf_rdat_b9c1_d3 };
  assign _0332_ = { cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41], cbuf_rd_sel_ram_d3[41:40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40], cbuf_rd_sel_ram_d3[40] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5535" *) { cbuf_rdat_b10c0_d3, cbuf_rdat_b10c1_d3 };
  assign _0333_ = { cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39], cbuf_rd_sel_ram_d3[39:38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38], cbuf_rd_sel_ram_d3[38] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5536" *) { cbuf_rdat_b11c0_d3, cbuf_rdat_b11c1_d3 };
  assign _0334_ = { cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37], cbuf_rd_sel_ram_d3[37:36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36], cbuf_rd_sel_ram_d3[36] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5537" *) { cbuf_rdat_b12c0_d3, cbuf_rdat_b12c1_d3 };
  assign _0335_ = { cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35], cbuf_rd_sel_ram_d3[35:34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34], cbuf_rd_sel_ram_d3[34] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5538" *) { cbuf_rdat_b13c0_d3, cbuf_rdat_b13c1_d3 };
  assign _0336_ = { cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33], cbuf_rd_sel_ram_d3[33:32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32], cbuf_rd_sel_ram_d3[32] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5539" *) { cbuf_rdat_b14c0_d3, cbuf_rdat_b14c1_d3 };
  assign _0337_ = { cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31], cbuf_rd_sel_ram_d3[31:30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30], cbuf_rd_sel_ram_d3[30] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5603" *) { cbuf_rdat_b1c0_d3, cbuf_rdat_b1c1_d3 };
  assign _0338_ = { cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29], cbuf_rd_sel_ram_d3[29:28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28], cbuf_rd_sel_ram_d3[28] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5604" *) { cbuf_rdat_b2c0_d3, cbuf_rdat_b2c1_d3 };
  assign _0339_ = { cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27], cbuf_rd_sel_ram_d3[27:26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26], cbuf_rd_sel_ram_d3[26] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5605" *) { cbuf_rdat_b3c0_d3, cbuf_rdat_b3c1_d3 };
  assign _0340_ = { cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25], cbuf_rd_sel_ram_d3[25:24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24], cbuf_rd_sel_ram_d3[24] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5606" *) { cbuf_rdat_b4c0_d3, cbuf_rdat_b4c1_d3 };
  assign _0341_ = { cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23], cbuf_rd_sel_ram_d3[23:22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22], cbuf_rd_sel_ram_d3[22] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5607" *) { cbuf_rdat_b5c0_d3, cbuf_rdat_b5c1_d3 };
  assign _0342_ = { cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21], cbuf_rd_sel_ram_d3[21:20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20], cbuf_rd_sel_ram_d3[20] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5608" *) { cbuf_rdat_b6c0_d3, cbuf_rdat_b6c1_d3 };
  assign _0343_ = { cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19], cbuf_rd_sel_ram_d3[19:18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18], cbuf_rd_sel_ram_d3[18] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5609" *) { cbuf_rdat_b7c0_d3, cbuf_rdat_b7c1_d3 };
  assign _0344_ = { cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17], cbuf_rd_sel_ram_d3[17:16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16], cbuf_rd_sel_ram_d3[16] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5610" *) { cbuf_rdat_b8c0_d3, cbuf_rdat_b8c1_d3 };
  assign _0345_ = { cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15], cbuf_rd_sel_ram_d3[15:14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14], cbuf_rd_sel_ram_d3[14] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5611" *) { cbuf_rdat_b9c0_d3, cbuf_rdat_b9c1_d3 };
  assign _0346_ = { cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13], cbuf_rd_sel_ram_d3[13:12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12], cbuf_rd_sel_ram_d3[12] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5612" *) { cbuf_rdat_b10c0_d3, cbuf_rdat_b10c1_d3 };
  assign _0347_ = { cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11], cbuf_rd_sel_ram_d3[11:10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10], cbuf_rd_sel_ram_d3[10] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5613" *) { cbuf_rdat_b11c0_d3, cbuf_rdat_b11c1_d3 };
  assign _0348_ = { cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9], cbuf_rd_sel_ram_d3[9:8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8], cbuf_rd_sel_ram_d3[8] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5614" *) { cbuf_rdat_b12c0_d3, cbuf_rdat_b12c1_d3 };
  assign _0349_ = { cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7], cbuf_rd_sel_ram_d3[7:6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6], cbuf_rd_sel_ram_d3[6] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5615" *) { cbuf_rdat_b13c0_d3, cbuf_rdat_b13c1_d3 };
  assign _0350_ = { cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5], cbuf_rd_sel_ram_d3[5:4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4], cbuf_rd_sel_ram_d3[4] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5616" *) { cbuf_rdat_b14c0_d3, cbuf_rdat_b14c1_d3 };
  assign _0351_ = { cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3], cbuf_rd_sel_ram_d3[3:2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2], cbuf_rd_sel_ram_d3[2] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5617" *) { cbuf_rdat_b15c0_d3, cbuf_rdat_b15c1_d3 };
  assign cbuf_p2_rd_data_d4_w = { cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1], cbuf_rd_sel_ram_d3[1:0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0], cbuf_rd_sel_ram_d3[0] } & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5625" *) { cbuf_rdat_b15c0_d3, cbuf_rdat_b15c1_d3 };
  assign cbuf_p0_wr_lo_en = cdma2buf_dat_wr_en & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:829" *) cdma2buf_dat_wr_hsel[0];
  assign cbuf_p0_wr_hi_en = cdma2buf_dat_wr_en & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:830" *) cdma2buf_dat_wr_hsel[1];
  assign cbuf_p1_wr_lo_en = cdma2buf_wt_wr_en & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:835" *) _0412_;
  assign cbuf_p1_wr_hi_en = cdma2buf_wt_wr_en & (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:836" *) cdma2buf_wt_wr_hsel;
  assign _0352_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1003" *) 4'b1010;
  assign _0353_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1010" *) 4'b1011;
  assign _0354_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1024" *) 4'b1100;
  assign _0355_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1038" *) 4'b1101;
  assign _0356_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1052" *) 4'b1110;
  assign _0357_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1066" *) 1'b1;
  assign _0358_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1080" *) 2'b10;
  assign _0359_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1094" *) 2'b11;
  assign _0360_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1108" *) 3'b100;
  assign _0361_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1122" *) 3'b101;
  assign _0362_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1136" *) 3'b110;
  assign _0363_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1150" *) 3'b111;
  assign _0364_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1164" *) 4'b1000;
  assign _0365_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1178" *) 4'b1001;
  assign _0366_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1192" *) 4'b1010;
  assign _0367_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1206" *) 4'b1011;
  assign _0368_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1220" *) 4'b1100;
  assign _0369_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1234" *) 4'b1101;
  assign _0370_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1248" *) 4'b1110;
  assign _0371_ = cdma2buf_wt_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1262" *) 4'b1111;
  assign _0372_ = ! (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3292" *) sc2buf_dat_rd_addr[11:8];
  assign _0373_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3306" *) 1'b1;
  assign _0374_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3320" *) 2'b10;
  assign _0375_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3334" *) 2'b11;
  assign _0376_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3348" *) 3'b100;
  assign _0377_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3362" *) 3'b101;
  assign _0378_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3376" *) 3'b110;
  assign _0379_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3390" *) 3'b111;
  assign _0380_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3404" *) 4'b1000;
  assign _0381_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3418" *) 4'b1001;
  assign _0382_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3432" *) 4'b1010;
  assign _0383_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3446" *) 4'b1011;
  assign _0384_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3460" *) 4'b1100;
  assign _0385_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3474" *) 4'b1101;
  assign _0386_ = sc2buf_dat_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3488" *) 4'b1110;
  assign _0387_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3502" *) 1'b1;
  assign _0388_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3516" *) 2'b10;
  assign _0389_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3530" *) 2'b11;
  assign _0390_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3544" *) 3'b100;
  assign _0391_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3558" *) 3'b101;
  assign _0392_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3572" *) 3'b110;
  assign _0393_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3586" *) 3'b111;
  assign _0394_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3600" *) 4'b1000;
  assign _0395_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3614" *) 4'b1001;
  assign _0396_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3628" *) 4'b1010;
  assign _0397_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3642" *) 4'b1011;
  assign _0398_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3656" *) 4'b1100;
  assign _0399_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3670" *) 4'b1101;
  assign _0400_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3684" *) 4'b1110;
  assign _0401_ = sc2buf_wt_rd_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3698" *) 4'b1111;
  assign _0402_ = ! (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:856" *) cdma2buf_dat_wr_addr[11:8];
  assign _0403_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:870" *) 1'b1;
  assign _0404_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:884" *) 2'b10;
  assign _0405_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:898" *) 2'b11;
  assign _0406_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:912" *) 3'b100;
  assign _0407_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:926" *) 3'b101;
  assign _0408_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:940" *) 3'b110;
  assign _0409_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:954" *) 3'b111;
  assign _0410_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:968" *) 4'b1000;
  assign _0411_ = cdma2buf_dat_wr_addr[11:8] == (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:982" *) 4'b1001;
  assign cbuf_p0_wr_sel_ram_b10c1_w = _0352_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1004" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b11c0_w = _0353_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1011" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b11c1_w = _0353_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1018" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b12c0_w = _0354_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1025" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b12c1_w = _0354_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1032" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b13c0_w = _0355_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1039" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b13c1_w = _0355_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1046" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b14c0_w = _0356_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1053" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b14c1_w = _0356_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1060" *) cbuf_p0_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b1c0_w = _0357_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1067" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b1c1_w = _0357_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1074" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b2c0_w = _0358_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1081" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b2c1_w = _0358_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1088" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b3c0_w = _0359_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1095" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b3c1_w = _0359_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1102" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b4c0_w = _0360_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1109" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b4c1_w = _0360_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1116" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b5c0_w = _0361_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1123" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b5c1_w = _0361_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1130" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b6c0_w = _0362_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1137" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b6c1_w = _0362_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1144" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b7c0_w = _0363_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1151" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b7c1_w = _0363_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1158" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b8c0_w = _0364_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1165" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b8c1_w = _0364_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1172" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b9c0_w = _0365_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1179" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b9c1_w = _0365_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1186" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b10c0_w = _0366_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1193" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b10c1_w = _0366_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1200" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b11c0_w = _0367_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1207" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b11c1_w = _0367_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1214" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b12c0_w = _0368_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1221" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b12c1_w = _0368_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1228" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b13c0_w = _0369_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1235" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b13c1_w = _0369_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1242" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b14c0_w = _0370_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1249" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b14c1_w = _0370_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1256" *) cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_sel_ram_b15c0_w = _0371_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1263" *) cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b15c1_w = _0371_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1270" *) cbuf_p1_wr_hi_en;
  assign cbuf_p0_rd_sel_ram_b0c0_w = _0372_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3293" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b1c0_w = _0373_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3307" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b2c0_w = _0374_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3321" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b3c0_w = _0375_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3335" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b4c0_w = _0376_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3349" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b5c0_w = _0377_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3363" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b6c0_w = _0378_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3377" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b7c0_w = _0379_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3391" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b8c0_w = _0380_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3405" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b9c0_w = _0381_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3419" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b10c0_w = _0382_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3433" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b11c0_w = _0383_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3447" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b12c0_w = _0384_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3461" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b13c0_w = _0385_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3475" *) sc2buf_dat_rd_en;
  assign cbuf_p0_rd_sel_ram_b14c0_w = _0386_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3489" *) sc2buf_dat_rd_en;
  assign cbuf_p1_rd_sel_ram_b1c0_w = _0387_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3503" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b2c0_w = _0388_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3517" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b3c0_w = _0389_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3531" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b4c0_w = _0390_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3545" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b5c0_w = _0391_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3559" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b6c0_w = _0392_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3573" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b7c0_w = _0393_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3587" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b8c0_w = _0394_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3601" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b9c0_w = _0395_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3615" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b10c0_w = _0396_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3629" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b11c0_w = _0397_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3643" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b12c0_w = _0398_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3657" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b13c0_w = _0399_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3671" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b14c0_w = _0400_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3685" *) sc2buf_wt_rd_en;
  assign cbuf_p1_rd_sel_ram_b15c0_w = _0401_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3699" *) sc2buf_wt_rd_en;
  assign cbuf_p0_wr_sel_ram_b0c0_w = _0402_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:857" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b0c1_w = _0402_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:864" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b1c0_w = _0403_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:871" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b1c1_w = _0403_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:878" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b2c0_w = _0404_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:885" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b2c1_w = _0404_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:892" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b3c0_w = _0405_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:899" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b3c1_w = _0405_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:906" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b4c0_w = _0406_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:913" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b4c1_w = _0406_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:920" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b5c0_w = _0407_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:927" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b5c1_w = _0407_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:934" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b6c0_w = _0408_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:941" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b6c1_w = _0408_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:948" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b7c0_w = _0409_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:955" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b7c1_w = _0409_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:962" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b8c0_w = _0410_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:969" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b8c1_w = _0410_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:976" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b9c0_w = _0411_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:983" *) cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b9c1_w = _0411_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:990" *) cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_sel_ram_b10c0_w = _0352_ && (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:997" *) cbuf_p0_wr_lo_en;
  assign _0412_ = ~ (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:835" *) cdma2buf_wt_wr_hsel;
  assign _0162_ = cbuf_p0_wr_sel_ram_b1c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1359" *) cbuf_p1_wr_sel_ram_b1c0_w;
  assign _0163_ = cbuf_p0_wr_sel_ram_b1c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1366" *) cbuf_p1_wr_sel_ram_b1c1_w;
  assign _0164_ = cbuf_p0_wr_sel_ram_b2c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1373" *) cbuf_p1_wr_sel_ram_b2c0_w;
  assign _0165_ = cbuf_p0_wr_sel_ram_b2c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1380" *) cbuf_p1_wr_sel_ram_b2c1_w;
  assign _0166_ = cbuf_p0_wr_sel_ram_b3c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1387" *) cbuf_p1_wr_sel_ram_b3c0_w;
  assign _0167_ = cbuf_p0_wr_sel_ram_b3c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1394" *) cbuf_p1_wr_sel_ram_b3c1_w;
  assign _0168_ = cbuf_p0_wr_sel_ram_b4c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1401" *) cbuf_p1_wr_sel_ram_b4c0_w;
  assign _0169_ = cbuf_p0_wr_sel_ram_b4c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1408" *) cbuf_p1_wr_sel_ram_b4c1_w;
  assign _0170_ = cbuf_p0_wr_sel_ram_b5c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1415" *) cbuf_p1_wr_sel_ram_b5c0_w;
  assign _0171_ = cbuf_p0_wr_sel_ram_b5c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1422" *) cbuf_p1_wr_sel_ram_b5c1_w;
  assign _0172_ = cbuf_p0_wr_sel_ram_b6c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1429" *) cbuf_p1_wr_sel_ram_b6c0_w;
  assign _0173_ = cbuf_p0_wr_sel_ram_b6c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1436" *) cbuf_p1_wr_sel_ram_b6c1_w;
  assign _0174_ = cbuf_p0_wr_sel_ram_b7c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1443" *) cbuf_p1_wr_sel_ram_b7c0_w;
  assign _0175_ = cbuf_p0_wr_sel_ram_b7c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1450" *) cbuf_p1_wr_sel_ram_b7c1_w;
  assign _0176_ = cbuf_p0_wr_sel_ram_b8c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1457" *) cbuf_p1_wr_sel_ram_b8c0_w;
  assign _0177_ = cbuf_p0_wr_sel_ram_b8c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1464" *) cbuf_p1_wr_sel_ram_b8c1_w;
  assign _0178_ = cbuf_p0_wr_sel_ram_b9c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1471" *) cbuf_p1_wr_sel_ram_b9c0_w;
  assign _0179_ = cbuf_p0_wr_sel_ram_b9c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1478" *) cbuf_p1_wr_sel_ram_b9c1_w;
  assign _0152_ = cbuf_p0_wr_sel_ram_b10c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1485" *) cbuf_p1_wr_sel_ram_b10c0_w;
  assign _0153_ = cbuf_p0_wr_sel_ram_b10c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1492" *) cbuf_p1_wr_sel_ram_b10c1_w;
  assign _0154_ = cbuf_p0_wr_sel_ram_b11c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1499" *) cbuf_p1_wr_sel_ram_b11c0_w;
  assign _0155_ = cbuf_p0_wr_sel_ram_b11c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1506" *) cbuf_p1_wr_sel_ram_b11c1_w;
  assign _0156_ = cbuf_p0_wr_sel_ram_b12c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1513" *) cbuf_p1_wr_sel_ram_b12c0_w;
  assign _0157_ = cbuf_p0_wr_sel_ram_b12c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1520" *) cbuf_p1_wr_sel_ram_b12c1_w;
  assign _0158_ = cbuf_p0_wr_sel_ram_b13c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1527" *) cbuf_p1_wr_sel_ram_b13c0_w;
  assign _0159_ = cbuf_p0_wr_sel_ram_b13c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1534" *) cbuf_p1_wr_sel_ram_b13c1_w;
  assign _0160_ = cbuf_p0_wr_sel_ram_b14c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1541" *) cbuf_p1_wr_sel_ram_b14c0_w;
  assign _0161_ = cbuf_p0_wr_sel_ram_b14c1_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1548" *) cbuf_p1_wr_sel_ram_b14c1_w;
  assign cbuf_wa_b1c0 = _0180_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1713" *) _0181_;
  assign cbuf_wdat_b1c0 = _0182_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1715" *) _0183_;
  assign cbuf_wa_b1c1 = _0184_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1726" *) _0185_;
  assign cbuf_wdat_b1c1 = _0186_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1728" *) _0187_;
  assign cbuf_wa_b2c0 = _0188_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1739" *) _0189_;
  assign cbuf_wdat_b2c0 = _0190_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1741" *) _0191_;
  assign cbuf_wa_b2c1 = _0192_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1752" *) _0193_;
  assign cbuf_wdat_b2c1 = _0194_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1754" *) _0195_;
  assign cbuf_wa_b3c0 = _0196_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1765" *) _0197_;
  assign cbuf_wdat_b3c0 = _0198_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1767" *) _0199_;
  assign cbuf_wa_b3c1 = _0200_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1778" *) _0201_;
  assign cbuf_wdat_b3c1 = _0202_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1780" *) _0203_;
  assign cbuf_wa_b4c0 = _0204_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1791" *) _0205_;
  assign cbuf_wdat_b4c0 = _0206_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1793" *) _0207_;
  assign cbuf_wa_b4c1 = _0208_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1804" *) _0209_;
  assign cbuf_wdat_b4c1 = _0210_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1806" *) _0211_;
  assign cbuf_wa_b5c0 = _0212_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1817" *) _0213_;
  assign cbuf_wdat_b5c0 = _0214_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1819" *) _0215_;
  assign cbuf_wa_b5c1 = _0216_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1830" *) _0217_;
  assign cbuf_wdat_b5c1 = _0218_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1832" *) _0219_;
  assign cbuf_wa_b6c0 = _0220_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1843" *) _0221_;
  assign cbuf_wdat_b6c0 = _0222_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1845" *) _0223_;
  assign cbuf_wa_b6c1 = _0224_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1856" *) _0225_;
  assign cbuf_wdat_b6c1 = _0226_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1858" *) _0227_;
  assign cbuf_wa_b7c0 = _0228_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1869" *) _0229_;
  assign cbuf_wdat_b7c0 = _0230_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1871" *) _0231_;
  assign cbuf_wa_b7c1 = _0232_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1882" *) _0233_;
  assign cbuf_wdat_b7c1 = _0234_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1884" *) _0235_;
  assign cbuf_wa_b8c0 = _0236_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1895" *) _0237_;
  assign cbuf_wdat_b8c0 = _0238_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1897" *) _0239_;
  assign cbuf_wa_b8c1 = _0240_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1908" *) _0241_;
  assign cbuf_wdat_b8c1 = _0242_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1910" *) _0243_;
  assign cbuf_wa_b9c0 = _0244_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1921" *) _0245_;
  assign cbuf_wdat_b9c0 = _0246_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1923" *) _0247_;
  assign cbuf_wa_b9c1 = _0248_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1934" *) _0249_;
  assign cbuf_wdat_b9c1 = _0250_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1936" *) _0251_;
  assign cbuf_wa_b10c0 = _0252_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1947" *) _0253_;
  assign cbuf_wdat_b10c0 = _0254_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1949" *) _0255_;
  assign cbuf_wa_b10c1 = _0256_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1960" *) _0257_;
  assign cbuf_wdat_b10c1 = _0258_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1962" *) _0259_;
  assign cbuf_wa_b11c0 = _0260_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1973" *) _0261_;
  assign cbuf_wdat_b11c0 = _0262_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1975" *) _0263_;
  assign cbuf_wa_b11c1 = _0264_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1986" *) _0265_;
  assign cbuf_wdat_b11c1 = _0266_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1988" *) _0267_;
  assign cbuf_wa_b12c0 = _0268_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1999" *) _0269_;
  assign cbuf_wdat_b12c0 = _0270_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2001" *) _0271_;
  assign cbuf_wa_b12c1 = _0272_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2012" *) _0273_;
  assign cbuf_wdat_b12c1 = _0274_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2014" *) _0275_;
  assign cbuf_wa_b13c0 = _0276_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2025" *) _0277_;
  assign cbuf_wdat_b13c0 = _0278_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2027" *) _0279_;
  assign cbuf_wa_b13c1 = _0280_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2038" *) _0281_;
  assign cbuf_wdat_b13c1 = _0282_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2040" *) _0283_;
  assign cbuf_wa_b14c0 = _0284_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2051" *) _0285_;
  assign cbuf_wdat_b14c0 = _0286_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2053" *) _0287_;
  assign cbuf_wa_b14c1 = _0288_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2064" *) _0289_;
  assign cbuf_wdat_b14c1 = _0290_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2066" *) _0291_;
  assign cbuf_re_b1c0_w = cbuf_p0_rd_sel_ram_b1c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3732" *) cbuf_p1_rd_sel_ram_b1c0_w;
  assign cbuf_re_b2c0_w = cbuf_p0_rd_sel_ram_b2c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3744" *) cbuf_p1_rd_sel_ram_b2c0_w;
  assign cbuf_re_b3c0_w = cbuf_p0_rd_sel_ram_b3c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3756" *) cbuf_p1_rd_sel_ram_b3c0_w;
  assign cbuf_re_b4c0_w = cbuf_p0_rd_sel_ram_b4c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3768" *) cbuf_p1_rd_sel_ram_b4c0_w;
  assign cbuf_re_b5c0_w = cbuf_p0_rd_sel_ram_b5c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3780" *) cbuf_p1_rd_sel_ram_b5c0_w;
  assign cbuf_re_b6c0_w = cbuf_p0_rd_sel_ram_b6c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3792" *) cbuf_p1_rd_sel_ram_b6c0_w;
  assign cbuf_re_b7c0_w = cbuf_p0_rd_sel_ram_b7c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3804" *) cbuf_p1_rd_sel_ram_b7c0_w;
  assign cbuf_re_b8c0_w = cbuf_p0_rd_sel_ram_b8c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3816" *) cbuf_p1_rd_sel_ram_b8c0_w;
  assign cbuf_re_b9c0_w = cbuf_p0_rd_sel_ram_b9c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3828" *) cbuf_p1_rd_sel_ram_b9c0_w;
  assign cbuf_re_b10c0_w = cbuf_p0_rd_sel_ram_b10c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3840" *) cbuf_p1_rd_sel_ram_b10c0_w;
  assign cbuf_re_b11c0_w = cbuf_p0_rd_sel_ram_b11c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3852" *) cbuf_p1_rd_sel_ram_b11c0_w;
  assign cbuf_re_b12c0_w = cbuf_p0_rd_sel_ram_b12c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3864" *) cbuf_p1_rd_sel_ram_b12c0_w;
  assign cbuf_re_b13c0_w = cbuf_p0_rd_sel_ram_b13c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3876" *) cbuf_p1_rd_sel_ram_b13c0_w;
  assign cbuf_re_b14c0_w = cbuf_p0_rd_sel_ram_b14c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3888" *) cbuf_p1_rd_sel_ram_b14c0_w;
  assign cbuf_re_b15c0_w = cbuf_p1_rd_sel_ram_b15c0_w | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3900" *) sc2buf_wmb_rd_en;
  assign cbuf_ra_b1c0_w = _0292_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3927" *) _0293_;
  assign cbuf_ra_b2c0_w = _0294_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3945" *) _0295_;
  assign cbuf_ra_b3c0_w = _0296_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3963" *) _0297_;
  assign cbuf_ra_b4c0_w = _0298_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3981" *) _0299_;
  assign cbuf_ra_b5c0_w = _0300_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3999" *) _0301_;
  assign cbuf_ra_b6c0_w = _0302_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4017" *) _0303_;
  assign cbuf_ra_b7c0_w = _0304_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4035" *) _0305_;
  assign cbuf_ra_b8c0_w = _0306_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4053" *) _0307_;
  assign cbuf_ra_b9c0_w = _0308_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4071" *) _0309_;
  assign cbuf_ra_b10c0_w = _0310_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4089" *) _0311_;
  assign cbuf_ra_b11c0_w = _0312_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4107" *) _0313_;
  assign cbuf_ra_b12c0_w = _0314_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4125" *) _0315_;
  assign cbuf_ra_b13c0_w = _0316_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4143" *) _0317_;
  assign cbuf_ra_b14c0_w = _0318_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4161" *) _0319_;
  assign cbuf_ra_b15c0_w = _0320_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4179" *) _0321_;
  assign _0413_ = _0322_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5526" *) _0323_;
  assign _0414_ = _0413_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5527" *) _0324_;
  assign _0415_ = _0414_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5528" *) _0325_;
  assign _0416_ = _0415_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5529" *) _0326_;
  assign _0417_ = _0416_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5530" *) _0327_;
  assign _0418_ = _0417_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5531" *) _0328_;
  assign _0419_ = _0418_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5532" *) _0329_;
  assign _0420_ = _0419_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5533" *) _0330_;
  assign _0421_ = _0420_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5534" *) _0331_;
  assign _0422_ = _0421_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5535" *) _0332_;
  assign _0423_ = _0422_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5536" *) _0333_;
  assign _0424_ = _0423_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5537" *) _0334_;
  assign _0425_ = _0424_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5538" *) _0335_;
  assign cbuf_p0_rd_data_d4_w = _0425_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5539" *) _0336_;
  assign _0426_ = _0337_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5604" *) _0338_;
  assign _0427_ = _0426_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5605" *) _0339_;
  assign _0428_ = _0427_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5606" *) _0340_;
  assign _0429_ = _0428_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5607" *) _0341_;
  assign _0430_ = _0429_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5608" *) _0342_;
  assign _0431_ = _0430_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5609" *) _0343_;
  assign _0432_ = _0431_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5610" *) _0344_;
  assign _0433_ = _0432_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5611" *) _0345_;
  assign _0434_ = _0433_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5612" *) _0346_;
  assign _0435_ = _0434_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5613" *) _0347_;
  assign _0436_ = _0435_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5614" *) _0348_;
  assign _0437_ = _0436_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5615" *) _0349_;
  assign _0438_ = _0437_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5616" *) _0350_;
  assign cbuf_p1_rd_data_d4_w = _0438_ | (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5617" *) _0351_;
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_data_d6[511:0] <= _0023_;
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_data_d6[1023:512] <= _0022_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_data_d6[511:0] <= _0014_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_data_d6[1023:512] <= _0013_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_data_d6[511:0] <= _0005_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_data_d6[1023:512] <= _0004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p2_rd_valid_d6 <= 1'b0;
    else
      cbuf_p2_rd_valid_d6 <= cbuf_p2_rd_en_d5;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p2_rd_en_d5 <= 1'b0;
    else
      cbuf_p2_rd_en_d5 <= cbuf_rd_en_d4[0];
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p1_rd_valid_d6 <= 1'b0;
    else
      cbuf_p1_rd_valid_d6 <= cbuf_p1_rd_en_d5;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p1_rd_en_d5 <= 1'b0;
    else
      cbuf_p1_rd_en_d5 <= cbuf_rd_en_d4[1];
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p0_rd_valid_d6 <= 1'b0;
    else
      cbuf_p0_rd_valid_d6 <= cbuf_p0_rd_en_d5;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_p0_rd_en_d5 <= 1'b0;
    else
      cbuf_p0_rd_en_d5 <= cbuf_rd_en_d4[2];
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_c1_data_d5 <= _0019_;
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_c0_data_d5 <= _0018_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_c1_data_d5 <= _0010_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_c0_data_d5 <= _0009_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_c1_data_d5 <= _0001_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_c0_data_d5 <= _0000_;
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_data_d4[1023:512] <= _0020_;
  always @(posedge nvdla_core_clk)
      cbuf_p2_rd_data_d4[511:0] <= _0021_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_data_d4[1023:512] <= _0011_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_rd_data_d4[511:0] <= _0012_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_data_d4[1023:512] <= _0002_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_rd_data_d4[511:0] <= _0003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_rd_en_d4 <= 3'b000;
    else
      cbuf_rd_en_d4 <= cbuf_rd_en_d3;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b15c1_d3 <= _0069_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b15c0_d3 <= _0068_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b14c1_d3 <= _0067_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b14c0_d3 <= _0066_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b13c1_d3 <= _0065_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b13c0_d3 <= _0064_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b12c1_d3 <= _0063_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b12c0_d3 <= _0062_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b11c1_d3 <= _0061_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b11c0_d3 <= _0060_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b10c1_d3 <= _0059_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b10c0_d3 <= _0058_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b9c1_d3 <= _0087_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b9c0_d3 <= _0086_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b8c1_d3 <= _0085_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b8c0_d3 <= _0084_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b7c1_d3 <= _0083_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b7c0_d3 <= _0082_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b6c1_d3 <= _0081_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b6c0_d3 <= _0080_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b5c1_d3 <= _0079_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b5c0_d3 <= _0078_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b4c1_d3 <= _0077_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b4c0_d3 <= _0076_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b3c1_d3 <= _0075_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b3c0_d3 <= _0074_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b2c1_d3 <= _0073_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b2c0_d3 <= _0072_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b1c1_d3 <= _0071_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b1c0_d3 <= _0070_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b0c1_d3 <= _0057_;
  always @(posedge nvdla_core_clk)
      cbuf_rdat_b0c0_d3 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_rd_en_d3 <= 3'b000;
    else
      cbuf_rd_en_d3 <= cbuf_rd_en_d2;
  reg [60:0] _0976_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      _0976_ <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    else
      _0976_ <= cbuf_rd_sel_ram_d2[60:0];
  assign cbuf_rd_sel_ram_d3[60:0] = _0976_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b15c1_d2 <= 1'b0;
    else
      cbuf_re_b15c1_d2 <= cbuf_re_b15c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b14c1_d2 <= 1'b0;
    else
      cbuf_re_b14c1_d2 <= cbuf_re_b14c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b13c1_d2 <= 1'b0;
    else
      cbuf_re_b13c1_d2 <= cbuf_re_b13c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b12c1_d2 <= 1'b0;
    else
      cbuf_re_b12c1_d2 <= cbuf_re_b12c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b11c1_d2 <= 1'b0;
    else
      cbuf_re_b11c1_d2 <= cbuf_re_b11c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b10c1_d2 <= 1'b0;
    else
      cbuf_re_b10c1_d2 <= cbuf_re_b10c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b9c1_d2 <= 1'b0;
    else
      cbuf_re_b9c1_d2 <= cbuf_re_b9c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b8c1_d2 <= 1'b0;
    else
      cbuf_re_b8c1_d2 <= cbuf_re_b8c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b7c1_d2 <= 1'b0;
    else
      cbuf_re_b7c1_d2 <= cbuf_re_b7c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b6c1_d2 <= 1'b0;
    else
      cbuf_re_b6c1_d2 <= cbuf_re_b6c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b5c1_d2 <= 1'b0;
    else
      cbuf_re_b5c1_d2 <= cbuf_re_b5c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b4c1_d2 <= 1'b0;
    else
      cbuf_re_b4c1_d2 <= cbuf_re_b4c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b3c1_d2 <= 1'b0;
    else
      cbuf_re_b3c1_d2 <= cbuf_re_b3c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b2c1_d2 <= 1'b0;
    else
      cbuf_re_b2c1_d2 <= cbuf_re_b2c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b1c1_d2 <= 1'b0;
    else
      cbuf_re_b1c1_d2 <= cbuf_re_b1c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b0c1_d2 <= 1'b0;
    else
      cbuf_re_b0c1_d2 <= cbuf_re_b0c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_rd_en_d2 <= 3'b000;
    else
      cbuf_rd_en_d2 <= cbuf_rd_en_d1;
  reg [60:0] _0994_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      _0994_ <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    else
      _0994_ <= cbuf_rd_sel_ram_d1[60:0];
  assign cbuf_rd_sel_ram_d2[60:0] = _0994_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b15c1 <= _0037_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b15c0 <= _0036_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b14c1 <= _0035_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b14c0 <= _0034_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b13c1 <= _0033_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b13c0 <= _0032_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b12c1 <= _0031_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b12c0 <= _0030_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b11c1 <= _0029_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b11c0 <= _0028_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b10c1 <= _0027_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b10c0 <= _0026_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b9c1 <= _0055_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b9c0 <= _0054_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b8c1 <= _0053_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b8c0 <= _0052_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b7c1 <= _0051_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b7c0 <= _0050_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b6c1 <= _0049_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b6c0 <= _0048_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b5c1 <= _0047_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b5c0 <= _0046_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b4c1 <= _0045_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b4c0 <= _0044_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b3c1 <= _0043_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b3c0 <= _0042_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b2c1 <= _0041_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b2c0 <= _0040_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b1c1 <= _0039_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b1c0 <= _0038_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b0c1 <= _0025_;
  always @(posedge nvdla_core_clk)
      cbuf_ra_b0c0 <= _0024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b15c1 <= 1'b0;
    else
      cbuf_re_b15c1 <= cbuf_re_b15c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b14c1 <= 1'b0;
    else
      cbuf_re_b14c1 <= cbuf_re_b14c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b13c1 <= 1'b0;
    else
      cbuf_re_b13c1 <= cbuf_re_b13c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b12c1 <= 1'b0;
    else
      cbuf_re_b12c1 <= cbuf_re_b12c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b11c1 <= 1'b0;
    else
      cbuf_re_b11c1 <= cbuf_re_b11c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b10c1 <= 1'b0;
    else
      cbuf_re_b10c1 <= cbuf_re_b10c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b9c1 <= 1'b0;
    else
      cbuf_re_b9c1 <= cbuf_re_b9c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b8c1 <= 1'b0;
    else
      cbuf_re_b8c1 <= cbuf_re_b8c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b7c1 <= 1'b0;
    else
      cbuf_re_b7c1 <= cbuf_re_b7c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b6c1 <= 1'b0;
    else
      cbuf_re_b6c1 <= cbuf_re_b6c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b5c1 <= 1'b0;
    else
      cbuf_re_b5c1 <= cbuf_re_b5c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b4c1 <= 1'b0;
    else
      cbuf_re_b4c1 <= cbuf_re_b4c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b3c1 <= 1'b0;
    else
      cbuf_re_b3c1 <= cbuf_re_b3c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b2c1 <= 1'b0;
    else
      cbuf_re_b2c1 <= cbuf_re_b2c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b1c1 <= 1'b0;
    else
      cbuf_re_b1c1 <= cbuf_re_b1c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_re_b0c1 <= 1'b0;
    else
      cbuf_re_b0c1 <= cbuf_p0_rd_sel_ram_b0c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_rd_en_d1 <= 3'b000;
    else
      cbuf_rd_en_d1 <= { sc2buf_dat_rd_en, sc2buf_wt_rd_en, sc2buf_wmb_rd_en };
  reg [60:0] _1044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      _1044_ <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    else
      _1044_ <= { cbuf_p0_rd_sel_ram_b0c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b1c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b2c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b3c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b4c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b5c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b6c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b7c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b8c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b9c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b10c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b11c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b12c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b13c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p0_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b1c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b2c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b3c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b4c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b5c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b6c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b7c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b8c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b9c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b10c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b11c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b12c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b13c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b14c0_w, cbuf_p1_rd_sel_ram_b15c0_w, cbuf_p1_rd_sel_ram_b15c0_w, sc2buf_wmb_rd_en, sc2buf_wmb_rd_en };
  assign cbuf_rd_sel_ram_d1[60:0] = _1044_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b15c1_d2 <= _0133_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b15c0_d2 <= _0132_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b14c1_d2 <= _0131_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b14c0_d2 <= _0130_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b13c1_d2 <= _0129_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b13c0_d2 <= _0128_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b12c1_d2 <= _0127_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b12c0_d2 <= _0126_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b11c1_d2 <= _0125_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b11c0_d2 <= _0124_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b10c1_d2 <= _0123_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b10c0_d2 <= _0122_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b9c1_d2 <= _0151_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b9c0_d2 <= _0150_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b8c1_d2 <= _0149_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b8c0_d2 <= _0148_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b7c1_d2 <= _0147_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b7c0_d2 <= _0146_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b6c1_d2 <= _0145_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b6c0_d2 <= _0144_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b5c1_d2 <= _0143_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b5c0_d2 <= _0142_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b4c1_d2 <= _0141_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b4c0_d2 <= _0140_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b3c1_d2 <= _0139_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b3c0_d2 <= _0138_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b2c1_d2 <= _0137_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b2c0_d2 <= _0136_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b1c1_d2 <= _0135_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b1c0_d2 <= _0134_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b0c1_d2 <= _0121_;
  always @(posedge nvdla_core_clk)
      cbuf_wdat_b0c0_d2 <= _0120_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b15c1_d2 <= _0101_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b15c0_d2 <= _0100_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b14c1_d2 <= _0099_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b14c0_d2 <= _0098_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b13c1_d2 <= _0097_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b13c0_d2 <= _0096_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b12c1_d2 <= _0095_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b12c0_d2 <= _0094_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b11c1_d2 <= _0093_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b11c0_d2 <= _0092_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b10c1_d2 <= _0091_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b10c0_d2 <= _0090_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b9c1_d2 <= _0119_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b9c0_d2 <= _0118_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b8c1_d2 <= _0117_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b8c0_d2 <= _0116_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b7c1_d2 <= _0115_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b7c0_d2 <= _0114_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b6c1_d2 <= _0113_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b6c0_d2 <= _0112_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b5c1_d2 <= _0111_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b5c0_d2 <= _0110_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b4c1_d2 <= _0109_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b4c0_d2 <= _0108_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b3c1_d2 <= _0107_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b3c0_d2 <= _0106_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b2c1_d2 <= _0105_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b2c0_d2 <= _0104_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b1c1_d2 <= _0103_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b1c0_d2 <= _0102_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b0c1_d2 <= _0089_;
  always @(posedge nvdla_core_clk)
      cbuf_wa_b0c0_d2 <= _0088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b15c1_d2 <= 1'b0;
    else
      cbuf_we_b15c1_d2 <= cbuf_we_b15c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b15c0_d2 <= 1'b0;
    else
      cbuf_we_b15c0_d2 <= cbuf_we_b15c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b14c1_d2 <= 1'b0;
    else
      cbuf_we_b14c1_d2 <= cbuf_we_b14c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b14c0_d2 <= 1'b0;
    else
      cbuf_we_b14c0_d2 <= cbuf_we_b14c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b13c1_d2 <= 1'b0;
    else
      cbuf_we_b13c1_d2 <= cbuf_we_b13c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b13c0_d2 <= 1'b0;
    else
      cbuf_we_b13c0_d2 <= cbuf_we_b13c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b12c1_d2 <= 1'b0;
    else
      cbuf_we_b12c1_d2 <= cbuf_we_b12c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b12c0_d2 <= 1'b0;
    else
      cbuf_we_b12c0_d2 <= cbuf_we_b12c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b11c1_d2 <= 1'b0;
    else
      cbuf_we_b11c1_d2 <= cbuf_we_b11c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b11c0_d2 <= 1'b0;
    else
      cbuf_we_b11c0_d2 <= cbuf_we_b11c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b10c1_d2 <= 1'b0;
    else
      cbuf_we_b10c1_d2 <= cbuf_we_b10c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b10c0_d2 <= 1'b0;
    else
      cbuf_we_b10c0_d2 <= cbuf_we_b10c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b9c1_d2 <= 1'b0;
    else
      cbuf_we_b9c1_d2 <= cbuf_we_b9c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b9c0_d2 <= 1'b0;
    else
      cbuf_we_b9c0_d2 <= cbuf_we_b9c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b8c1_d2 <= 1'b0;
    else
      cbuf_we_b8c1_d2 <= cbuf_we_b8c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b8c0_d2 <= 1'b0;
    else
      cbuf_we_b8c0_d2 <= cbuf_we_b8c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b7c1_d2 <= 1'b0;
    else
      cbuf_we_b7c1_d2 <= cbuf_we_b7c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b7c0_d2 <= 1'b0;
    else
      cbuf_we_b7c0_d2 <= cbuf_we_b7c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b6c1_d2 <= 1'b0;
    else
      cbuf_we_b6c1_d2 <= cbuf_we_b6c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b6c0_d2 <= 1'b0;
    else
      cbuf_we_b6c0_d2 <= cbuf_we_b6c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b5c1_d2 <= 1'b0;
    else
      cbuf_we_b5c1_d2 <= cbuf_we_b5c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b5c0_d2 <= 1'b0;
    else
      cbuf_we_b5c0_d2 <= cbuf_we_b5c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b4c1_d2 <= 1'b0;
    else
      cbuf_we_b4c1_d2 <= cbuf_we_b4c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b4c0_d2 <= 1'b0;
    else
      cbuf_we_b4c0_d2 <= cbuf_we_b4c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b3c1_d2 <= 1'b0;
    else
      cbuf_we_b3c1_d2 <= cbuf_we_b3c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b3c0_d2 <= 1'b0;
    else
      cbuf_we_b3c0_d2 <= cbuf_we_b3c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b2c1_d2 <= 1'b0;
    else
      cbuf_we_b2c1_d2 <= cbuf_we_b2c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b2c0_d2 <= 1'b0;
    else
      cbuf_we_b2c0_d2 <= cbuf_we_b2c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b1c1_d2 <= 1'b0;
    else
      cbuf_we_b1c1_d2 <= cbuf_we_b1c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b1c0_d2 <= 1'b0;
    else
      cbuf_we_b1c0_d2 <= cbuf_we_b1c0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b0c1_d2 <= 1'b0;
    else
      cbuf_we_b0c1_d2 <= cbuf_we_b0c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b0c0_d2 <= 1'b0;
    else
      cbuf_we_b0c0_d2 <= cbuf_we_b0c0;
  always @(posedge nvdla_core_clk)
      cbuf_p1_wr_hi_data_d1 <= _0016_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_wr_lo_data_d1 <= _0017_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_wr_hi_data_d1 <= _0007_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_wr_lo_data_d1 <= _0008_;
  always @(posedge nvdla_core_clk)
      cbuf_p1_wr_addr_d1 <= _0015_;
  always @(posedge nvdla_core_clk)
      cbuf_p0_wr_addr_d1 <= _0006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b15c1 <= 1'b0;
    else
      cbuf_we_b15c1 <= cbuf_p1_wr_sel_ram_b15c1_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b15c0 <= 1'b0;
    else
      cbuf_we_b15c0 <= cbuf_p1_wr_sel_ram_b15c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b14c1 <= 1'b0;
    else
      cbuf_we_b14c1 <= _0161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b14c0 <= 1'b0;
    else
      cbuf_we_b14c0 <= _0160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b13c1 <= 1'b0;
    else
      cbuf_we_b13c1 <= _0159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b13c0 <= 1'b0;
    else
      cbuf_we_b13c0 <= _0158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b12c1 <= 1'b0;
    else
      cbuf_we_b12c1 <= _0157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b12c0 <= 1'b0;
    else
      cbuf_we_b12c0 <= _0156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b11c1 <= 1'b0;
    else
      cbuf_we_b11c1 <= _0155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b11c0 <= 1'b0;
    else
      cbuf_we_b11c0 <= _0154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b10c1 <= 1'b0;
    else
      cbuf_we_b10c1 <= _0153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b10c0 <= 1'b0;
    else
      cbuf_we_b10c0 <= _0152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b9c1 <= 1'b0;
    else
      cbuf_we_b9c1 <= _0179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b9c0 <= 1'b0;
    else
      cbuf_we_b9c0 <= _0178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b8c1 <= 1'b0;
    else
      cbuf_we_b8c1 <= _0177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b8c0 <= 1'b0;
    else
      cbuf_we_b8c0 <= _0176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b7c1 <= 1'b0;
    else
      cbuf_we_b7c1 <= _0175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b7c0 <= 1'b0;
    else
      cbuf_we_b7c0 <= _0174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b6c1 <= 1'b0;
    else
      cbuf_we_b6c1 <= _0173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b6c0 <= 1'b0;
    else
      cbuf_we_b6c0 <= _0172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b5c1 <= 1'b0;
    else
      cbuf_we_b5c1 <= _0171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b5c0 <= 1'b0;
    else
      cbuf_we_b5c0 <= _0170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b4c1 <= 1'b0;
    else
      cbuf_we_b4c1 <= _0169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b4c0 <= 1'b0;
    else
      cbuf_we_b4c0 <= _0168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b3c1 <= 1'b0;
    else
      cbuf_we_b3c1 <= _0167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b3c0 <= 1'b0;
    else
      cbuf_we_b3c0 <= _0166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b2c1 <= 1'b0;
    else
      cbuf_we_b2c1 <= _0165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b2c0 <= 1'b0;
    else
      cbuf_we_b2c0 <= _0164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b1c1 <= 1'b0;
    else
      cbuf_we_b1c1 <= _0163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b1c0 <= 1'b0;
    else
      cbuf_we_b1c0 <= _0162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b0c1 <= 1'b0;
    else
      cbuf_we_b0c1 <= cbuf_p0_wr_sel_ram_b0c1_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_we_b0c0 <= 1'b0;
    else
      cbuf_we_b0c0 <= cbuf_p0_wr_sel_ram_b0c0_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cbuf_wr_sel_ram_d1 <= 60'b000000000000000000000000000000000000000000000000000000000000;
    else
      cbuf_wr_sel_ram_d1 <= { cbuf_p0_wr_sel_ram_b0c0_w, cbuf_p0_wr_sel_ram_b0c1_w, cbuf_p0_wr_sel_ram_b1c0_w, cbuf_p0_wr_sel_ram_b1c1_w, cbuf_p0_wr_sel_ram_b2c0_w, cbuf_p0_wr_sel_ram_b2c1_w, cbuf_p0_wr_sel_ram_b3c0_w, cbuf_p0_wr_sel_ram_b3c1_w, cbuf_p0_wr_sel_ram_b4c0_w, cbuf_p0_wr_sel_ram_b4c1_w, cbuf_p0_wr_sel_ram_b5c0_w, cbuf_p0_wr_sel_ram_b5c1_w, cbuf_p0_wr_sel_ram_b6c0_w, cbuf_p0_wr_sel_ram_b6c1_w, cbuf_p0_wr_sel_ram_b7c0_w, cbuf_p0_wr_sel_ram_b7c1_w, cbuf_p0_wr_sel_ram_b8c0_w, cbuf_p0_wr_sel_ram_b8c1_w, cbuf_p0_wr_sel_ram_b9c0_w, cbuf_p0_wr_sel_ram_b9c1_w, cbuf_p0_wr_sel_ram_b10c0_w, cbuf_p0_wr_sel_ram_b10c1_w, cbuf_p0_wr_sel_ram_b11c0_w, cbuf_p0_wr_sel_ram_b11c1_w, cbuf_p0_wr_sel_ram_b12c0_w, cbuf_p0_wr_sel_ram_b12c1_w, cbuf_p0_wr_sel_ram_b13c0_w, cbuf_p0_wr_sel_ram_b13c1_w, cbuf_p0_wr_sel_ram_b14c0_w, cbuf_p0_wr_sel_ram_b14c1_w, cbuf_p1_wr_sel_ram_b1c0_w, cbuf_p1_wr_sel_ram_b1c1_w, cbuf_p1_wr_sel_ram_b2c0_w, cbuf_p1_wr_sel_ram_b2c1_w, cbuf_p1_wr_sel_ram_b3c0_w, cbuf_p1_wr_sel_ram_b3c1_w, cbuf_p1_wr_sel_ram_b4c0_w, cbuf_p1_wr_sel_ram_b4c1_w, cbuf_p1_wr_sel_ram_b5c0_w, cbuf_p1_wr_sel_ram_b5c1_w, cbuf_p1_wr_sel_ram_b6c0_w, cbuf_p1_wr_sel_ram_b6c1_w, cbuf_p1_wr_sel_ram_b7c0_w, cbuf_p1_wr_sel_ram_b7c1_w, cbuf_p1_wr_sel_ram_b8c0_w, cbuf_p1_wr_sel_ram_b8c1_w, cbuf_p1_wr_sel_ram_b9c0_w, cbuf_p1_wr_sel_ram_b9c1_w, cbuf_p1_wr_sel_ram_b10c0_w, cbuf_p1_wr_sel_ram_b10c1_w, cbuf_p1_wr_sel_ram_b11c0_w, cbuf_p1_wr_sel_ram_b11c1_w, cbuf_p1_wr_sel_ram_b12c0_w, cbuf_p1_wr_sel_ram_b12c1_w, cbuf_p1_wr_sel_ram_b13c0_w, cbuf_p1_wr_sel_ram_b13c1_w, cbuf_p1_wr_sel_ram_b14c0_w, cbuf_p1_wr_sel_ram_b14c1_w, cbuf_p1_wr_sel_ram_b15c0_w, cbuf_p1_wr_sel_ram_b15c1_w };
  assign _0023_ = cbuf_p2_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5897" *) cbuf_p2_rd_c0_data_d5 : cbuf_p2_rd_data_d6[511:0];
  assign _0022_ = cbuf_p2_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5892" *) cbuf_p2_rd_c1_data_d5 : cbuf_p2_rd_data_d6[1023:512];
  assign _0014_ = cbuf_p1_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5887" *) cbuf_p1_rd_c0_data_d5 : cbuf_p1_rd_data_d6[511:0];
  assign _0013_ = cbuf_p1_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5882" *) cbuf_p1_rd_c1_data_d5 : cbuf_p1_rd_data_d6[1023:512];
  assign _0005_ = cbuf_p0_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5877" *) cbuf_p0_rd_c0_data_d5 : cbuf_p0_rd_data_d6[511:0];
  assign _0004_ = cbuf_p0_rd_en_d5 ? (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5872" *) cbuf_p0_rd_c1_data_d5 : cbuf_p0_rd_data_d6[1023:512];
  assign _0019_ = cbuf_rd_en_d4[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5815" *) cbuf_p2_rd_data_d4[511:0] : cbuf_p2_rd_c1_data_d5;
  assign _0018_ = cbuf_rd_en_d4[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5796" *) cbuf_p2_rd_data_d4[1023:512] : cbuf_p2_rd_c0_data_d5;
  assign _0010_ = cbuf_rd_en_d4[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5777" *) cbuf_p1_rd_data_d4[511:0] : cbuf_p1_rd_c1_data_d5;
  assign _0009_ = cbuf_rd_en_d4[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5758" *) cbuf_p1_rd_data_d4[1023:512] : cbuf_p1_rd_c0_data_d5;
  assign _0001_ = cbuf_rd_en_d4[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5739" *) cbuf_p0_rd_data_d4[511:0] : cbuf_p0_rd_c1_data_d5;
  assign _0000_ = cbuf_rd_en_d4[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5720" *) cbuf_p0_rd_data_d4[1023:512] : cbuf_p0_rd_c0_data_d5;
  assign _0020_ = cbuf_rd_en_d3[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5688" *) cbuf_p2_rd_data_d4_w[1023:512] : cbuf_p2_rd_data_d4[1023:512];
  assign _0021_ = cbuf_rd_en_d3[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5678" *) cbuf_p2_rd_data_d4_w[511:0] : cbuf_p2_rd_data_d4[511:0];
  assign _0011_ = cbuf_rd_en_d3[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5668" *) cbuf_p1_rd_data_d4_w[1023:512] : cbuf_p1_rd_data_d4[1023:512];
  assign _0012_ = cbuf_rd_en_d3[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5658" *) cbuf_p1_rd_data_d4_w[511:0] : cbuf_p1_rd_data_d4[511:0];
  assign _0002_ = cbuf_rd_en_d3[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5648" *) cbuf_p0_rd_data_d4_w[1023:512] : cbuf_p0_rd_data_d4[1023:512];
  assign _0003_ = cbuf_rd_en_d3[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5638" *) cbuf_p0_rd_data_d4_w[511:0] : cbuf_p0_rd_data_d4[511:0];
  assign _0069_ = cbuf_re_b15c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5386" *) cbuf_rdat_b15c1 : cbuf_rdat_b15c1_d3;
  assign _0068_ = cbuf_re_b15c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5376" *) cbuf_rdat_b15c0 : cbuf_rdat_b15c0_d3;
  assign _0067_ = cbuf_re_b14c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5366" *) cbuf_rdat_b14c1 : cbuf_rdat_b14c1_d3;
  assign _0066_ = cbuf_re_b14c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5356" *) cbuf_rdat_b14c0 : cbuf_rdat_b14c0_d3;
  assign _0065_ = cbuf_re_b13c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5346" *) cbuf_rdat_b13c1 : cbuf_rdat_b13c1_d3;
  assign _0064_ = cbuf_re_b13c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5336" *) cbuf_rdat_b13c0 : cbuf_rdat_b13c0_d3;
  assign _0063_ = cbuf_re_b12c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5326" *) cbuf_rdat_b12c1 : cbuf_rdat_b12c1_d3;
  assign _0062_ = cbuf_re_b12c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5316" *) cbuf_rdat_b12c0 : cbuf_rdat_b12c0_d3;
  assign _0061_ = cbuf_re_b11c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5306" *) cbuf_rdat_b11c1 : cbuf_rdat_b11c1_d3;
  assign _0060_ = cbuf_re_b11c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5296" *) cbuf_rdat_b11c0 : cbuf_rdat_b11c0_d3;
  assign _0059_ = cbuf_re_b10c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5286" *) cbuf_rdat_b10c1 : cbuf_rdat_b10c1_d3;
  assign _0058_ = cbuf_re_b10c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5276" *) cbuf_rdat_b10c0 : cbuf_rdat_b10c0_d3;
  assign _0087_ = cbuf_re_b9c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5266" *) cbuf_rdat_b9c1 : cbuf_rdat_b9c1_d3;
  assign _0086_ = cbuf_re_b9c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5256" *) cbuf_rdat_b9c0 : cbuf_rdat_b9c0_d3;
  assign _0085_ = cbuf_re_b8c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5246" *) cbuf_rdat_b8c1 : cbuf_rdat_b8c1_d3;
  assign _0084_ = cbuf_re_b8c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5236" *) cbuf_rdat_b8c0 : cbuf_rdat_b8c0_d3;
  assign _0083_ = cbuf_re_b7c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5226" *) cbuf_rdat_b7c1 : cbuf_rdat_b7c1_d3;
  assign _0082_ = cbuf_re_b7c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5216" *) cbuf_rdat_b7c0 : cbuf_rdat_b7c0_d3;
  assign _0081_ = cbuf_re_b6c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5206" *) cbuf_rdat_b6c1 : cbuf_rdat_b6c1_d3;
  assign _0080_ = cbuf_re_b6c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5196" *) cbuf_rdat_b6c0 : cbuf_rdat_b6c0_d3;
  assign _0079_ = cbuf_re_b5c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5186" *) cbuf_rdat_b5c1 : cbuf_rdat_b5c1_d3;
  assign _0078_ = cbuf_re_b5c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5176" *) cbuf_rdat_b5c0 : cbuf_rdat_b5c0_d3;
  assign _0077_ = cbuf_re_b4c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5166" *) cbuf_rdat_b4c1 : cbuf_rdat_b4c1_d3;
  assign _0076_ = cbuf_re_b4c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5156" *) cbuf_rdat_b4c0 : cbuf_rdat_b4c0_d3;
  assign _0075_ = cbuf_re_b3c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5146" *) cbuf_rdat_b3c1 : cbuf_rdat_b3c1_d3;
  assign _0074_ = cbuf_re_b3c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5136" *) cbuf_rdat_b3c0 : cbuf_rdat_b3c0_d3;
  assign _0073_ = cbuf_re_b2c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5126" *) cbuf_rdat_b2c1 : cbuf_rdat_b2c1_d3;
  assign _0072_ = cbuf_re_b2c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5116" *) cbuf_rdat_b2c0 : cbuf_rdat_b2c0_d3;
  assign _0071_ = cbuf_re_b1c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5106" *) cbuf_rdat_b1c1 : cbuf_rdat_b1c1_d3;
  assign _0070_ = cbuf_re_b1c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5096" *) cbuf_rdat_b1c0 : cbuf_rdat_b1c0_d3;
  assign _0057_ = cbuf_re_b0c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5086" *) cbuf_rdat_b0c1 : cbuf_rdat_b0c1_d3;
  assign _0056_ = cbuf_re_b0c1_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:5076" *) cbuf_rdat_b0c0 : cbuf_rdat_b0c0_d3;
  assign _0037_ = cbuf_re_b15c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4805" *) cbuf_ra_b15c0_w : cbuf_ra_b15c1;
  assign _0036_ = cbuf_re_b15c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4795" *) cbuf_ra_b15c0_w : cbuf_ra_b15c0;
  assign _0035_ = cbuf_re_b14c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4785" *) cbuf_ra_b14c0_w : cbuf_ra_b14c1;
  assign _0034_ = cbuf_re_b14c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4775" *) cbuf_ra_b14c0_w : cbuf_ra_b14c0;
  assign _0033_ = cbuf_re_b13c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4765" *) cbuf_ra_b13c0_w : cbuf_ra_b13c1;
  assign _0032_ = cbuf_re_b13c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4755" *) cbuf_ra_b13c0_w : cbuf_ra_b13c0;
  assign _0031_ = cbuf_re_b12c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4745" *) cbuf_ra_b12c0_w : cbuf_ra_b12c1;
  assign _0030_ = cbuf_re_b12c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4735" *) cbuf_ra_b12c0_w : cbuf_ra_b12c0;
  assign _0029_ = cbuf_re_b11c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4725" *) cbuf_ra_b11c0_w : cbuf_ra_b11c1;
  assign _0028_ = cbuf_re_b11c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4715" *) cbuf_ra_b11c0_w : cbuf_ra_b11c0;
  assign _0027_ = cbuf_re_b10c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4705" *) cbuf_ra_b10c0_w : cbuf_ra_b10c1;
  assign _0026_ = cbuf_re_b10c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4695" *) cbuf_ra_b10c0_w : cbuf_ra_b10c0;
  assign _0055_ = cbuf_re_b9c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4685" *) cbuf_ra_b9c0_w : cbuf_ra_b9c1;
  assign _0054_ = cbuf_re_b9c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4675" *) cbuf_ra_b9c0_w : cbuf_ra_b9c0;
  assign _0053_ = cbuf_re_b8c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4665" *) cbuf_ra_b8c0_w : cbuf_ra_b8c1;
  assign _0052_ = cbuf_re_b8c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4655" *) cbuf_ra_b8c0_w : cbuf_ra_b8c0;
  assign _0051_ = cbuf_re_b7c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4645" *) cbuf_ra_b7c0_w : cbuf_ra_b7c1;
  assign _0050_ = cbuf_re_b7c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4635" *) cbuf_ra_b7c0_w : cbuf_ra_b7c0;
  assign _0049_ = cbuf_re_b6c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4625" *) cbuf_ra_b6c0_w : cbuf_ra_b6c1;
  assign _0048_ = cbuf_re_b6c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4615" *) cbuf_ra_b6c0_w : cbuf_ra_b6c0;
  assign _0047_ = cbuf_re_b5c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4605" *) cbuf_ra_b5c0_w : cbuf_ra_b5c1;
  assign _0046_ = cbuf_re_b5c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4595" *) cbuf_ra_b5c0_w : cbuf_ra_b5c0;
  assign _0045_ = cbuf_re_b4c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4585" *) cbuf_ra_b4c0_w : cbuf_ra_b4c1;
  assign _0044_ = cbuf_re_b4c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4575" *) cbuf_ra_b4c0_w : cbuf_ra_b4c0;
  assign _0043_ = cbuf_re_b3c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4565" *) cbuf_ra_b3c0_w : cbuf_ra_b3c1;
  assign _0042_ = cbuf_re_b3c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4555" *) cbuf_ra_b3c0_w : cbuf_ra_b3c0;
  assign _0041_ = cbuf_re_b2c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4545" *) cbuf_ra_b2c0_w : cbuf_ra_b2c1;
  assign _0040_ = cbuf_re_b2c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4535" *) cbuf_ra_b2c0_w : cbuf_ra_b2c0;
  assign _0039_ = cbuf_re_b1c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4525" *) cbuf_ra_b1c0_w : cbuf_ra_b1c1;
  assign _0038_ = cbuf_re_b1c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4515" *) cbuf_ra_b1c0_w : cbuf_ra_b1c0;
  assign _0025_ = cbuf_p0_rd_sel_ram_b0c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4505" *) cbuf_ra_b0c0_w : cbuf_ra_b0c1;
  assign _0024_ = cbuf_p0_rd_sel_ram_b0c0_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:4495" *) cbuf_ra_b0c0_w : cbuf_ra_b0c0;
  assign _0133_ = cbuf_we_b15c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2942" *) cbuf_wdat_b15c1 : cbuf_wdat_b15c1_d2;
  assign _0132_ = cbuf_we_b15c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2932" *) cbuf_wdat_b15c0 : cbuf_wdat_b15c0_d2;
  assign _0131_ = cbuf_we_b14c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2922" *) cbuf_wdat_b14c1 : cbuf_wdat_b14c1_d2;
  assign _0130_ = cbuf_we_b14c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2912" *) cbuf_wdat_b14c0 : cbuf_wdat_b14c0_d2;
  assign _0129_ = cbuf_we_b13c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2902" *) cbuf_wdat_b13c1 : cbuf_wdat_b13c1_d2;
  assign _0128_ = cbuf_we_b13c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2892" *) cbuf_wdat_b13c0 : cbuf_wdat_b13c0_d2;
  assign _0127_ = cbuf_we_b12c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2882" *) cbuf_wdat_b12c1 : cbuf_wdat_b12c1_d2;
  assign _0126_ = cbuf_we_b12c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2872" *) cbuf_wdat_b12c0 : cbuf_wdat_b12c0_d2;
  assign _0125_ = cbuf_we_b11c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2862" *) cbuf_wdat_b11c1 : cbuf_wdat_b11c1_d2;
  assign _0124_ = cbuf_we_b11c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2852" *) cbuf_wdat_b11c0 : cbuf_wdat_b11c0_d2;
  assign _0123_ = cbuf_we_b10c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2842" *) cbuf_wdat_b10c1 : cbuf_wdat_b10c1_d2;
  assign _0122_ = cbuf_we_b10c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2832" *) cbuf_wdat_b10c0 : cbuf_wdat_b10c0_d2;
  assign _0151_ = cbuf_we_b9c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2822" *) cbuf_wdat_b9c1 : cbuf_wdat_b9c1_d2;
  assign _0150_ = cbuf_we_b9c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2812" *) cbuf_wdat_b9c0 : cbuf_wdat_b9c0_d2;
  assign _0149_ = cbuf_we_b8c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2802" *) cbuf_wdat_b8c1 : cbuf_wdat_b8c1_d2;
  assign _0148_ = cbuf_we_b8c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2792" *) cbuf_wdat_b8c0 : cbuf_wdat_b8c0_d2;
  assign _0147_ = cbuf_we_b7c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2782" *) cbuf_wdat_b7c1 : cbuf_wdat_b7c1_d2;
  assign _0146_ = cbuf_we_b7c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2772" *) cbuf_wdat_b7c0 : cbuf_wdat_b7c0_d2;
  assign _0145_ = cbuf_we_b6c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2762" *) cbuf_wdat_b6c1 : cbuf_wdat_b6c1_d2;
  assign _0144_ = cbuf_we_b6c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2752" *) cbuf_wdat_b6c0 : cbuf_wdat_b6c0_d2;
  assign _0143_ = cbuf_we_b5c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2742" *) cbuf_wdat_b5c1 : cbuf_wdat_b5c1_d2;
  assign _0142_ = cbuf_we_b5c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2732" *) cbuf_wdat_b5c0 : cbuf_wdat_b5c0_d2;
  assign _0141_ = cbuf_we_b4c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2722" *) cbuf_wdat_b4c1 : cbuf_wdat_b4c1_d2;
  assign _0140_ = cbuf_we_b4c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2712" *) cbuf_wdat_b4c0 : cbuf_wdat_b4c0_d2;
  assign _0139_ = cbuf_we_b3c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2702" *) cbuf_wdat_b3c1 : cbuf_wdat_b3c1_d2;
  assign _0138_ = cbuf_we_b3c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2692" *) cbuf_wdat_b3c0 : cbuf_wdat_b3c0_d2;
  assign _0137_ = cbuf_we_b2c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2682" *) cbuf_wdat_b2c1 : cbuf_wdat_b2c1_d2;
  assign _0136_ = cbuf_we_b2c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2672" *) cbuf_wdat_b2c0 : cbuf_wdat_b2c0_d2;
  assign _0135_ = cbuf_we_b1c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2662" *) cbuf_wdat_b1c1 : cbuf_wdat_b1c1_d2;
  assign _0134_ = cbuf_we_b1c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2652" *) cbuf_wdat_b1c0 : cbuf_wdat_b1c0_d2;
  assign _0121_ = cbuf_we_b0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2642" *) cbuf_wdat_b0c1 : cbuf_wdat_b0c1_d2;
  assign _0120_ = cbuf_we_b0c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2632" *) cbuf_wdat_b0c0 : cbuf_wdat_b0c0_d2;
  assign _0101_ = cbuf_we_b15c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2622" *) cbuf_wa_b15c1 : cbuf_wa_b15c1_d2;
  assign _0100_ = cbuf_we_b15c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2612" *) cbuf_wa_b15c0 : cbuf_wa_b15c0_d2;
  assign _0099_ = cbuf_we_b14c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2602" *) cbuf_wa_b14c1 : cbuf_wa_b14c1_d2;
  assign _0098_ = cbuf_we_b14c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2592" *) cbuf_wa_b14c0 : cbuf_wa_b14c0_d2;
  assign _0097_ = cbuf_we_b13c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2582" *) cbuf_wa_b13c1 : cbuf_wa_b13c1_d2;
  assign _0096_ = cbuf_we_b13c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2572" *) cbuf_wa_b13c0 : cbuf_wa_b13c0_d2;
  assign _0095_ = cbuf_we_b12c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2562" *) cbuf_wa_b12c1 : cbuf_wa_b12c1_d2;
  assign _0094_ = cbuf_we_b12c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2552" *) cbuf_wa_b12c0 : cbuf_wa_b12c0_d2;
  assign _0093_ = cbuf_we_b11c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2542" *) cbuf_wa_b11c1 : cbuf_wa_b11c1_d2;
  assign _0092_ = cbuf_we_b11c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2532" *) cbuf_wa_b11c0 : cbuf_wa_b11c0_d2;
  assign _0091_ = cbuf_we_b10c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2522" *) cbuf_wa_b10c1 : cbuf_wa_b10c1_d2;
  assign _0090_ = cbuf_we_b10c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2512" *) cbuf_wa_b10c0 : cbuf_wa_b10c0_d2;
  assign _0119_ = cbuf_we_b9c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2502" *) cbuf_wa_b9c1 : cbuf_wa_b9c1_d2;
  assign _0118_ = cbuf_we_b9c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2492" *) cbuf_wa_b9c0 : cbuf_wa_b9c0_d2;
  assign _0117_ = cbuf_we_b8c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2482" *) cbuf_wa_b8c1 : cbuf_wa_b8c1_d2;
  assign _0116_ = cbuf_we_b8c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2472" *) cbuf_wa_b8c0 : cbuf_wa_b8c0_d2;
  assign _0115_ = cbuf_we_b7c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2462" *) cbuf_wa_b7c1 : cbuf_wa_b7c1_d2;
  assign _0114_ = cbuf_we_b7c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2452" *) cbuf_wa_b7c0 : cbuf_wa_b7c0_d2;
  assign _0113_ = cbuf_we_b6c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2442" *) cbuf_wa_b6c1 : cbuf_wa_b6c1_d2;
  assign _0112_ = cbuf_we_b6c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2432" *) cbuf_wa_b6c0 : cbuf_wa_b6c0_d2;
  assign _0111_ = cbuf_we_b5c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2422" *) cbuf_wa_b5c1 : cbuf_wa_b5c1_d2;
  assign _0110_ = cbuf_we_b5c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2412" *) cbuf_wa_b5c0 : cbuf_wa_b5c0_d2;
  assign _0109_ = cbuf_we_b4c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2402" *) cbuf_wa_b4c1 : cbuf_wa_b4c1_d2;
  assign _0108_ = cbuf_we_b4c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2392" *) cbuf_wa_b4c0 : cbuf_wa_b4c0_d2;
  assign _0107_ = cbuf_we_b3c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2382" *) cbuf_wa_b3c1 : cbuf_wa_b3c1_d2;
  assign _0106_ = cbuf_we_b3c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2372" *) cbuf_wa_b3c0 : cbuf_wa_b3c0_d2;
  assign _0105_ = cbuf_we_b2c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2362" *) cbuf_wa_b2c1 : cbuf_wa_b2c1_d2;
  assign _0104_ = cbuf_we_b2c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2352" *) cbuf_wa_b2c0 : cbuf_wa_b2c0_d2;
  assign _0103_ = cbuf_we_b1c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2342" *) cbuf_wa_b1c1 : cbuf_wa_b1c1_d2;
  assign _0102_ = cbuf_we_b1c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2332" *) cbuf_wa_b1c0 : cbuf_wa_b1c0_d2;
  assign _0089_ = cbuf_we_b0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2322" *) cbuf_wa_b0c1 : cbuf_wa_b0c1_d2;
  assign _0088_ = cbuf_we_b0c0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2312" *) cbuf_wa_b0c0 : cbuf_wa_b0c0_d2;
  assign _0016_ = cbuf_p1_wr_hi_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1616" *) cdma2buf_wt_wr_data : cbuf_p1_wr_hi_data_d1;
  assign _0017_ = cbuf_p1_wr_lo_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1606" *) cdma2buf_wt_wr_data : cbuf_p1_wr_lo_data_d1;
  assign _0007_ = cbuf_p0_wr_hi_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1596" *) cdma2buf_dat_wr_data[1023:512] : cbuf_p0_wr_hi_data_d1;
  assign _0008_ = cbuf_p0_wr_lo_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1586" *) cdma2buf_dat_wr_data[511:0] : cbuf_p0_wr_lo_data_d1;
  assign _0015_ = cdma2buf_wt_wr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1576" *) cdma2buf_wt_wr_addr[7:0] : cbuf_p1_wr_addr_d1;
  assign _0006_ = cdma2buf_dat_wr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:1566" *) cdma2buf_dat_wr_addr[7:0] : cbuf_p0_wr_addr_d1;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2954" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank0_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b0c0_d2),
    .dout(cbuf_rdat_b0c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b0c0),
    .re(cbuf_re_b0c1),
    .wa(cbuf_wa_b0c0_d2),
    .we(cbuf_we_b0c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2964" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank0_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b0c1_d2),
    .dout(cbuf_rdat_b0c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b0c1),
    .re(cbuf_re_b0c1),
    .wa(cbuf_wa_b0c1_d2),
    .we(cbuf_we_b0c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3154" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank10_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b10c0_d2),
    .dout(cbuf_rdat_b10c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b10c0),
    .re(cbuf_re_b10c1),
    .wa(cbuf_wa_b10c0_d2),
    .we(cbuf_we_b10c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3164" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank10_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b10c1_d2),
    .dout(cbuf_rdat_b10c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b10c1),
    .re(cbuf_re_b10c1),
    .wa(cbuf_wa_b10c1_d2),
    .we(cbuf_we_b10c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3174" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank11_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b11c0_d2),
    .dout(cbuf_rdat_b11c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b11c0),
    .re(cbuf_re_b11c1),
    .wa(cbuf_wa_b11c0_d2),
    .we(cbuf_we_b11c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3184" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank11_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b11c1_d2),
    .dout(cbuf_rdat_b11c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b11c1),
    .re(cbuf_re_b11c1),
    .wa(cbuf_wa_b11c1_d2),
    .we(cbuf_we_b11c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3194" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank12_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b12c0_d2),
    .dout(cbuf_rdat_b12c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b12c0),
    .re(cbuf_re_b12c1),
    .wa(cbuf_wa_b12c0_d2),
    .we(cbuf_we_b12c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3204" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank12_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b12c1_d2),
    .dout(cbuf_rdat_b12c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b12c1),
    .re(cbuf_re_b12c1),
    .wa(cbuf_wa_b12c1_d2),
    .we(cbuf_we_b12c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3214" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank13_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b13c0_d2),
    .dout(cbuf_rdat_b13c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b13c0),
    .re(cbuf_re_b13c1),
    .wa(cbuf_wa_b13c0_d2),
    .we(cbuf_we_b13c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3224" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank13_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b13c1_d2),
    .dout(cbuf_rdat_b13c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b13c1),
    .re(cbuf_re_b13c1),
    .wa(cbuf_wa_b13c1_d2),
    .we(cbuf_we_b13c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3234" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank14_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b14c0_d2),
    .dout(cbuf_rdat_b14c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b14c0),
    .re(cbuf_re_b14c1),
    .wa(cbuf_wa_b14c0_d2),
    .we(cbuf_we_b14c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3244" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank14_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b14c1_d2),
    .dout(cbuf_rdat_b14c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b14c1),
    .re(cbuf_re_b14c1),
    .wa(cbuf_wa_b14c1_d2),
    .we(cbuf_we_b14c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3254" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank15_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b15c0_d2),
    .dout(cbuf_rdat_b15c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b15c0),
    .re(cbuf_re_b15c1),
    .wa(cbuf_wa_b15c0_d2),
    .we(cbuf_we_b15c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3264" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank15_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b15c1_d2),
    .dout(cbuf_rdat_b15c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b15c1),
    .re(cbuf_re_b15c1),
    .wa(cbuf_wa_b15c1_d2),
    .we(cbuf_we_b15c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2974" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank1_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b1c0_d2),
    .dout(cbuf_rdat_b1c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b1c0),
    .re(cbuf_re_b1c1),
    .wa(cbuf_wa_b1c0_d2),
    .we(cbuf_we_b1c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2984" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank1_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b1c1_d2),
    .dout(cbuf_rdat_b1c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b1c1),
    .re(cbuf_re_b1c1),
    .wa(cbuf_wa_b1c1_d2),
    .we(cbuf_we_b1c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:2994" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank2_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b2c0_d2),
    .dout(cbuf_rdat_b2c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b2c0),
    .re(cbuf_re_b2c1),
    .wa(cbuf_wa_b2c0_d2),
    .we(cbuf_we_b2c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3004" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank2_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b2c1_d2),
    .dout(cbuf_rdat_b2c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b2c1),
    .re(cbuf_re_b2c1),
    .wa(cbuf_wa_b2c1_d2),
    .we(cbuf_we_b2c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3014" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank3_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b3c0_d2),
    .dout(cbuf_rdat_b3c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b3c0),
    .re(cbuf_re_b3c1),
    .wa(cbuf_wa_b3c0_d2),
    .we(cbuf_we_b3c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3024" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank3_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b3c1_d2),
    .dout(cbuf_rdat_b3c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b3c1),
    .re(cbuf_re_b3c1),
    .wa(cbuf_wa_b3c1_d2),
    .we(cbuf_we_b3c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3034" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank4_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b4c0_d2),
    .dout(cbuf_rdat_b4c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b4c0),
    .re(cbuf_re_b4c1),
    .wa(cbuf_wa_b4c0_d2),
    .we(cbuf_we_b4c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3044" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank4_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b4c1_d2),
    .dout(cbuf_rdat_b4c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b4c1),
    .re(cbuf_re_b4c1),
    .wa(cbuf_wa_b4c1_d2),
    .we(cbuf_we_b4c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3054" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank5_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b5c0_d2),
    .dout(cbuf_rdat_b5c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b5c0),
    .re(cbuf_re_b5c1),
    .wa(cbuf_wa_b5c0_d2),
    .we(cbuf_we_b5c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3064" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank5_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b5c1_d2),
    .dout(cbuf_rdat_b5c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b5c1),
    .re(cbuf_re_b5c1),
    .wa(cbuf_wa_b5c1_d2),
    .we(cbuf_we_b5c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3074" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank6_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b6c0_d2),
    .dout(cbuf_rdat_b6c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b6c0),
    .re(cbuf_re_b6c1),
    .wa(cbuf_wa_b6c0_d2),
    .we(cbuf_we_b6c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3084" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank6_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b6c1_d2),
    .dout(cbuf_rdat_b6c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b6c1),
    .re(cbuf_re_b6c1),
    .wa(cbuf_wa_b6c1_d2),
    .we(cbuf_we_b6c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3094" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank7_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b7c0_d2),
    .dout(cbuf_rdat_b7c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b7c0),
    .re(cbuf_re_b7c1),
    .wa(cbuf_wa_b7c0_d2),
    .we(cbuf_we_b7c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3104" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank7_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b7c1_d2),
    .dout(cbuf_rdat_b7c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b7c1),
    .re(cbuf_re_b7c1),
    .wa(cbuf_wa_b7c1_d2),
    .we(cbuf_we_b7c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3114" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank8_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b8c0_d2),
    .dout(cbuf_rdat_b8c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b8c0),
    .re(cbuf_re_b8c1),
    .wa(cbuf_wa_b8c0_d2),
    .we(cbuf_we_b8c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3124" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank8_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b8c1_d2),
    .dout(cbuf_rdat_b8c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b8c1),
    .re(cbuf_re_b8c1),
    .wa(cbuf_wa_b8c1_d2),
    .we(cbuf_we_b8c1_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3134" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank9_column0 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b9c0_d2),
    .dout(cbuf_rdat_b9c0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b9c0),
    .re(cbuf_re_b9c1),
    .wa(cbuf_wa_b9c0_d2),
    .we(cbuf_we_b9c0_d2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cbuf/NV_NVDLA_cbuf.v:3144" *)
  nv_ram_rws_256x512 u_cbuf_ram_bank9_column1 (
    .clk(nvdla_core_clk),
    .di(cbuf_wdat_b9c1_d2),
    .dout(cbuf_rdat_b9c1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(cbuf_ra_b9c1),
    .re(cbuf_re_b9c1),
    .wa(cbuf_wa_b9c1_d2),
    .we(cbuf_we_b9c1_d2)
  );
  assign cbuf_p0_rd_addr = sc2buf_dat_rd_addr;
  assign cbuf_p0_rd_bank = sc2buf_dat_rd_addr[11:8];
  assign cbuf_p0_rd_c0_data_d4 = cbuf_p0_rd_data_d4[1023:512];
  assign cbuf_p0_rd_c0_data_d6_w = cbuf_p0_rd_c0_data_d5;
  assign cbuf_p0_rd_c0_valid_d5 = cbuf_p0_rd_en_d5;
  assign cbuf_p0_rd_c0_valid_d6_w = cbuf_p0_rd_en_d5;
  assign cbuf_p0_rd_c1_data_d4 = cbuf_p0_rd_data_d4[511:0];
  assign cbuf_p0_rd_c1_data_d6_w = cbuf_p0_rd_c1_data_d5;
  assign cbuf_p0_rd_c1_valid_d5 = cbuf_p0_rd_en_d5;
  assign cbuf_p0_rd_c1_valid_d6_w = cbuf_p0_rd_en_d5;
  assign cbuf_p0_rd_en = sc2buf_dat_rd_en;
  assign cbuf_p0_rd_en_d3 = cbuf_rd_en_d3[2];
  assign cbuf_p0_rd_en_d4 = cbuf_rd_en_d4[2];
  assign cbuf_p0_rd_sel_ram_b0c0_d3 = cbuf_rd_sel_ram_d3[60];
  assign cbuf_p0_rd_sel_ram_b0c1_d3 = cbuf_rd_sel_ram_d3[60];
  assign cbuf_p0_rd_sel_ram_b0c1_w = cbuf_p0_rd_sel_ram_b0c0_w;
  assign cbuf_p0_rd_sel_ram_b10c0_d3 = cbuf_rd_sel_ram_d3[41];
  assign cbuf_p0_rd_sel_ram_b10c1_d3 = cbuf_rd_sel_ram_d3[40];
  assign cbuf_p0_rd_sel_ram_b10c1_w = cbuf_p0_rd_sel_ram_b10c0_w;
  assign cbuf_p0_rd_sel_ram_b11c0_d3 = cbuf_rd_sel_ram_d3[39];
  assign cbuf_p0_rd_sel_ram_b11c1_d3 = cbuf_rd_sel_ram_d3[38];
  assign cbuf_p0_rd_sel_ram_b11c1_w = cbuf_p0_rd_sel_ram_b11c0_w;
  assign cbuf_p0_rd_sel_ram_b12c0_d3 = cbuf_rd_sel_ram_d3[37];
  assign cbuf_p0_rd_sel_ram_b12c1_d3 = cbuf_rd_sel_ram_d3[36];
  assign cbuf_p0_rd_sel_ram_b12c1_w = cbuf_p0_rd_sel_ram_b12c0_w;
  assign cbuf_p0_rd_sel_ram_b13c0_d3 = cbuf_rd_sel_ram_d3[35];
  assign cbuf_p0_rd_sel_ram_b13c1_d3 = cbuf_rd_sel_ram_d3[34];
  assign cbuf_p0_rd_sel_ram_b13c1_w = cbuf_p0_rd_sel_ram_b13c0_w;
  assign cbuf_p0_rd_sel_ram_b14c0_d3 = cbuf_rd_sel_ram_d3[33];
  assign cbuf_p0_rd_sel_ram_b14c1_d3 = cbuf_rd_sel_ram_d3[32];
  assign cbuf_p0_rd_sel_ram_b14c1_w = cbuf_p0_rd_sel_ram_b14c0_w;
  assign cbuf_p0_rd_sel_ram_b1c0_d3 = cbuf_rd_sel_ram_d3[59];
  assign cbuf_p0_rd_sel_ram_b1c1_d3 = cbuf_rd_sel_ram_d3[58];
  assign cbuf_p0_rd_sel_ram_b1c1_w = cbuf_p0_rd_sel_ram_b1c0_w;
  assign cbuf_p0_rd_sel_ram_b2c0_d3 = cbuf_rd_sel_ram_d3[57];
  assign cbuf_p0_rd_sel_ram_b2c1_d3 = cbuf_rd_sel_ram_d3[56];
  assign cbuf_p0_rd_sel_ram_b2c1_w = cbuf_p0_rd_sel_ram_b2c0_w;
  assign cbuf_p0_rd_sel_ram_b3c0_d3 = cbuf_rd_sel_ram_d3[55];
  assign cbuf_p0_rd_sel_ram_b3c1_d3 = cbuf_rd_sel_ram_d3[54];
  assign cbuf_p0_rd_sel_ram_b3c1_w = cbuf_p0_rd_sel_ram_b3c0_w;
  assign cbuf_p0_rd_sel_ram_b4c0_d3 = cbuf_rd_sel_ram_d3[53];
  assign cbuf_p0_rd_sel_ram_b4c1_d3 = cbuf_rd_sel_ram_d3[52];
  assign cbuf_p0_rd_sel_ram_b4c1_w = cbuf_p0_rd_sel_ram_b4c0_w;
  assign cbuf_p0_rd_sel_ram_b5c0_d3 = cbuf_rd_sel_ram_d3[51];
  assign cbuf_p0_rd_sel_ram_b5c1_d3 = cbuf_rd_sel_ram_d3[50];
  assign cbuf_p0_rd_sel_ram_b5c1_w = cbuf_p0_rd_sel_ram_b5c0_w;
  assign cbuf_p0_rd_sel_ram_b6c0_d3 = cbuf_rd_sel_ram_d3[49];
  assign cbuf_p0_rd_sel_ram_b6c1_d3 = cbuf_rd_sel_ram_d3[48];
  assign cbuf_p0_rd_sel_ram_b6c1_w = cbuf_p0_rd_sel_ram_b6c0_w;
  assign cbuf_p0_rd_sel_ram_b7c0_d3 = cbuf_rd_sel_ram_d3[47];
  assign cbuf_p0_rd_sel_ram_b7c1_d3 = cbuf_rd_sel_ram_d3[46];
  assign cbuf_p0_rd_sel_ram_b7c1_w = cbuf_p0_rd_sel_ram_b7c0_w;
  assign cbuf_p0_rd_sel_ram_b8c0_d3 = cbuf_rd_sel_ram_d3[45];
  assign cbuf_p0_rd_sel_ram_b8c1_d3 = cbuf_rd_sel_ram_d3[44];
  assign cbuf_p0_rd_sel_ram_b8c1_w = cbuf_p0_rd_sel_ram_b8c0_w;
  assign cbuf_p0_rd_sel_ram_b9c0_d3 = cbuf_rd_sel_ram_d3[43];
  assign cbuf_p0_rd_sel_ram_b9c1_d3 = cbuf_rd_sel_ram_d3[42];
  assign cbuf_p0_rd_sel_ram_b9c1_w = cbuf_p0_rd_sel_ram_b9c0_w;
  assign cbuf_p0_wr_addr = cdma2buf_dat_wr_addr;
  assign cbuf_p0_wr_bank = cdma2buf_dat_wr_addr[11:8];
  assign cbuf_p0_wr_en = cdma2buf_dat_wr_en;
  assign cbuf_p0_wr_hi_data = cdma2buf_dat_wr_data[1023:512];
  assign cbuf_p0_wr_hi_data_d1_w = cdma2buf_dat_wr_data[1023:512];
  assign cbuf_p0_wr_hi_en_d1_w = cbuf_p0_wr_hi_en;
  assign cbuf_p0_wr_lo_data = cdma2buf_dat_wr_data[511:0];
  assign cbuf_p0_wr_lo_data_d1_w = cdma2buf_dat_wr_data[511:0];
  assign cbuf_p0_wr_lo_en_d1_w = cbuf_p0_wr_lo_en;
  assign cbuf_p0_wr_sel_ram_b0c0_d1 = cbuf_wr_sel_ram_d1[59];
  assign cbuf_p0_wr_sel_ram_b0c1_d1 = cbuf_wr_sel_ram_d1[58];
  assign cbuf_p0_wr_sel_ram_b10c0_d1 = cbuf_wr_sel_ram_d1[39];
  assign cbuf_p0_wr_sel_ram_b10c1_d1 = cbuf_wr_sel_ram_d1[38];
  assign cbuf_p0_wr_sel_ram_b11c0_d1 = cbuf_wr_sel_ram_d1[37];
  assign cbuf_p0_wr_sel_ram_b11c1_d1 = cbuf_wr_sel_ram_d1[36];
  assign cbuf_p0_wr_sel_ram_b12c0_d1 = cbuf_wr_sel_ram_d1[35];
  assign cbuf_p0_wr_sel_ram_b12c1_d1 = cbuf_wr_sel_ram_d1[34];
  assign cbuf_p0_wr_sel_ram_b13c0_d1 = cbuf_wr_sel_ram_d1[33];
  assign cbuf_p0_wr_sel_ram_b13c1_d1 = cbuf_wr_sel_ram_d1[32];
  assign cbuf_p0_wr_sel_ram_b14c0_d1 = cbuf_wr_sel_ram_d1[31];
  assign cbuf_p0_wr_sel_ram_b14c1_d1 = cbuf_wr_sel_ram_d1[30];
  assign cbuf_p0_wr_sel_ram_b1c0_d1 = cbuf_wr_sel_ram_d1[57];
  assign cbuf_p0_wr_sel_ram_b1c1_d1 = cbuf_wr_sel_ram_d1[56];
  assign cbuf_p0_wr_sel_ram_b2c0_d1 = cbuf_wr_sel_ram_d1[55];
  assign cbuf_p0_wr_sel_ram_b2c1_d1 = cbuf_wr_sel_ram_d1[54];
  assign cbuf_p0_wr_sel_ram_b3c0_d1 = cbuf_wr_sel_ram_d1[53];
  assign cbuf_p0_wr_sel_ram_b3c1_d1 = cbuf_wr_sel_ram_d1[52];
  assign cbuf_p0_wr_sel_ram_b4c0_d1 = cbuf_wr_sel_ram_d1[51];
  assign cbuf_p0_wr_sel_ram_b4c1_d1 = cbuf_wr_sel_ram_d1[50];
  assign cbuf_p0_wr_sel_ram_b5c0_d1 = cbuf_wr_sel_ram_d1[49];
  assign cbuf_p0_wr_sel_ram_b5c1_d1 = cbuf_wr_sel_ram_d1[48];
  assign cbuf_p0_wr_sel_ram_b6c0_d1 = cbuf_wr_sel_ram_d1[47];
  assign cbuf_p0_wr_sel_ram_b6c1_d1 = cbuf_wr_sel_ram_d1[46];
  assign cbuf_p0_wr_sel_ram_b7c0_d1 = cbuf_wr_sel_ram_d1[45];
  assign cbuf_p0_wr_sel_ram_b7c1_d1 = cbuf_wr_sel_ram_d1[44];
  assign cbuf_p0_wr_sel_ram_b8c0_d1 = cbuf_wr_sel_ram_d1[43];
  assign cbuf_p0_wr_sel_ram_b8c1_d1 = cbuf_wr_sel_ram_d1[42];
  assign cbuf_p0_wr_sel_ram_b9c0_d1 = cbuf_wr_sel_ram_d1[41];
  assign cbuf_p0_wr_sel_ram_b9c1_d1 = cbuf_wr_sel_ram_d1[40];
  assign cbuf_p1_rd_addr = sc2buf_wt_rd_addr;
  assign cbuf_p1_rd_bank = sc2buf_wt_rd_addr[11:8];
  assign cbuf_p1_rd_c0_data_d4 = cbuf_p1_rd_data_d4[1023:512];
  assign cbuf_p1_rd_c0_data_d6_w = cbuf_p1_rd_c0_data_d5;
  assign cbuf_p1_rd_c0_valid_d5 = cbuf_p1_rd_en_d5;
  assign cbuf_p1_rd_c0_valid_d6_w = cbuf_p1_rd_en_d5;
  assign cbuf_p1_rd_c1_data_d4 = cbuf_p1_rd_data_d4[511:0];
  assign cbuf_p1_rd_c1_data_d6_w = cbuf_p1_rd_c1_data_d5;
  assign cbuf_p1_rd_c1_valid_d5 = cbuf_p1_rd_en_d5;
  assign cbuf_p1_rd_c1_valid_d6_w = cbuf_p1_rd_en_d5;
  assign cbuf_p1_rd_en = sc2buf_wt_rd_en;
  assign cbuf_p1_rd_en_d3 = cbuf_rd_en_d3[1];
  assign cbuf_p1_rd_en_d4 = cbuf_rd_en_d4[1];
  assign cbuf_p1_rd_sel_ram_b10c0_d3 = cbuf_rd_sel_ram_d3[13];
  assign cbuf_p1_rd_sel_ram_b10c1_d3 = cbuf_rd_sel_ram_d3[12];
  assign cbuf_p1_rd_sel_ram_b10c1_w = cbuf_p1_rd_sel_ram_b10c0_w;
  assign cbuf_p1_rd_sel_ram_b11c0_d3 = cbuf_rd_sel_ram_d3[11];
  assign cbuf_p1_rd_sel_ram_b11c1_d3 = cbuf_rd_sel_ram_d3[10];
  assign cbuf_p1_rd_sel_ram_b11c1_w = cbuf_p1_rd_sel_ram_b11c0_w;
  assign cbuf_p1_rd_sel_ram_b12c0_d3 = cbuf_rd_sel_ram_d3[9];
  assign cbuf_p1_rd_sel_ram_b12c1_d3 = cbuf_rd_sel_ram_d3[8];
  assign cbuf_p1_rd_sel_ram_b12c1_w = cbuf_p1_rd_sel_ram_b12c0_w;
  assign cbuf_p1_rd_sel_ram_b13c0_d3 = cbuf_rd_sel_ram_d3[7];
  assign cbuf_p1_rd_sel_ram_b13c1_d3 = cbuf_rd_sel_ram_d3[6];
  assign cbuf_p1_rd_sel_ram_b13c1_w = cbuf_p1_rd_sel_ram_b13c0_w;
  assign cbuf_p1_rd_sel_ram_b14c0_d3 = cbuf_rd_sel_ram_d3[5];
  assign cbuf_p1_rd_sel_ram_b14c1_d3 = cbuf_rd_sel_ram_d3[4];
  assign cbuf_p1_rd_sel_ram_b14c1_w = cbuf_p1_rd_sel_ram_b14c0_w;
  assign cbuf_p1_rd_sel_ram_b15c0_d3 = cbuf_rd_sel_ram_d3[3];
  assign cbuf_p1_rd_sel_ram_b15c1_d3 = cbuf_rd_sel_ram_d3[2];
  assign cbuf_p1_rd_sel_ram_b15c1_w = cbuf_p1_rd_sel_ram_b15c0_w;
  assign cbuf_p1_rd_sel_ram_b1c0_d3 = cbuf_rd_sel_ram_d3[31];
  assign cbuf_p1_rd_sel_ram_b1c1_d3 = cbuf_rd_sel_ram_d3[30];
  assign cbuf_p1_rd_sel_ram_b1c1_w = cbuf_p1_rd_sel_ram_b1c0_w;
  assign cbuf_p1_rd_sel_ram_b2c0_d3 = cbuf_rd_sel_ram_d3[29];
  assign cbuf_p1_rd_sel_ram_b2c1_d3 = cbuf_rd_sel_ram_d3[28];
  assign cbuf_p1_rd_sel_ram_b2c1_w = cbuf_p1_rd_sel_ram_b2c0_w;
  assign cbuf_p1_rd_sel_ram_b3c0_d3 = cbuf_rd_sel_ram_d3[27];
  assign cbuf_p1_rd_sel_ram_b3c1_d3 = cbuf_rd_sel_ram_d3[26];
  assign cbuf_p1_rd_sel_ram_b3c1_w = cbuf_p1_rd_sel_ram_b3c0_w;
  assign cbuf_p1_rd_sel_ram_b4c0_d3 = cbuf_rd_sel_ram_d3[25];
  assign cbuf_p1_rd_sel_ram_b4c1_d3 = cbuf_rd_sel_ram_d3[24];
  assign cbuf_p1_rd_sel_ram_b4c1_w = cbuf_p1_rd_sel_ram_b4c0_w;
  assign cbuf_p1_rd_sel_ram_b5c0_d3 = cbuf_rd_sel_ram_d3[23];
  assign cbuf_p1_rd_sel_ram_b5c1_d3 = cbuf_rd_sel_ram_d3[22];
  assign cbuf_p1_rd_sel_ram_b5c1_w = cbuf_p1_rd_sel_ram_b5c0_w;
  assign cbuf_p1_rd_sel_ram_b6c0_d3 = cbuf_rd_sel_ram_d3[21];
  assign cbuf_p1_rd_sel_ram_b6c1_d3 = cbuf_rd_sel_ram_d3[20];
  assign cbuf_p1_rd_sel_ram_b6c1_w = cbuf_p1_rd_sel_ram_b6c0_w;
  assign cbuf_p1_rd_sel_ram_b7c0_d3 = cbuf_rd_sel_ram_d3[19];
  assign cbuf_p1_rd_sel_ram_b7c1_d3 = cbuf_rd_sel_ram_d3[18];
  assign cbuf_p1_rd_sel_ram_b7c1_w = cbuf_p1_rd_sel_ram_b7c0_w;
  assign cbuf_p1_rd_sel_ram_b8c0_d3 = cbuf_rd_sel_ram_d3[17];
  assign cbuf_p1_rd_sel_ram_b8c1_d3 = cbuf_rd_sel_ram_d3[16];
  assign cbuf_p1_rd_sel_ram_b8c1_w = cbuf_p1_rd_sel_ram_b8c0_w;
  assign cbuf_p1_rd_sel_ram_b9c0_d3 = cbuf_rd_sel_ram_d3[15];
  assign cbuf_p1_rd_sel_ram_b9c1_d3 = cbuf_rd_sel_ram_d3[14];
  assign cbuf_p1_rd_sel_ram_b9c1_w = cbuf_p1_rd_sel_ram_b9c0_w;
  assign cbuf_p1_wr_addr = cdma2buf_wt_wr_addr;
  assign cbuf_p1_wr_bank = cdma2buf_wt_wr_addr[11:8];
  assign cbuf_p1_wr_data = cdma2buf_wt_wr_data;
  assign cbuf_p1_wr_en = cdma2buf_wt_wr_en;
  assign cbuf_p1_wr_hi_data_d1_w = cdma2buf_wt_wr_data;
  assign cbuf_p1_wr_hi_en_d1_w = cbuf_p1_wr_hi_en;
  assign cbuf_p1_wr_lo_data_d1_w = cdma2buf_wt_wr_data;
  assign cbuf_p1_wr_lo_en_d1_w = cbuf_p1_wr_lo_en;
  assign cbuf_p1_wr_sel_ram_b10c0_d1 = cbuf_wr_sel_ram_d1[11];
  assign cbuf_p1_wr_sel_ram_b10c1_d1 = cbuf_wr_sel_ram_d1[10];
  assign cbuf_p1_wr_sel_ram_b11c0_d1 = cbuf_wr_sel_ram_d1[9];
  assign cbuf_p1_wr_sel_ram_b11c1_d1 = cbuf_wr_sel_ram_d1[8];
  assign cbuf_p1_wr_sel_ram_b12c0_d1 = cbuf_wr_sel_ram_d1[7];
  assign cbuf_p1_wr_sel_ram_b12c1_d1 = cbuf_wr_sel_ram_d1[6];
  assign cbuf_p1_wr_sel_ram_b13c0_d1 = cbuf_wr_sel_ram_d1[5];
  assign cbuf_p1_wr_sel_ram_b13c1_d1 = cbuf_wr_sel_ram_d1[4];
  assign cbuf_p1_wr_sel_ram_b14c0_d1 = cbuf_wr_sel_ram_d1[3];
  assign cbuf_p1_wr_sel_ram_b14c1_d1 = cbuf_wr_sel_ram_d1[2];
  assign cbuf_p1_wr_sel_ram_b15c0_d1 = cbuf_wr_sel_ram_d1[1];
  assign cbuf_p1_wr_sel_ram_b15c1_d1 = cbuf_wr_sel_ram_d1[0];
  assign cbuf_p1_wr_sel_ram_b1c0_d1 = cbuf_wr_sel_ram_d1[29];
  assign cbuf_p1_wr_sel_ram_b1c1_d1 = cbuf_wr_sel_ram_d1[28];
  assign cbuf_p1_wr_sel_ram_b2c0_d1 = cbuf_wr_sel_ram_d1[27];
  assign cbuf_p1_wr_sel_ram_b2c1_d1 = cbuf_wr_sel_ram_d1[26];
  assign cbuf_p1_wr_sel_ram_b3c0_d1 = cbuf_wr_sel_ram_d1[25];
  assign cbuf_p1_wr_sel_ram_b3c1_d1 = cbuf_wr_sel_ram_d1[24];
  assign cbuf_p1_wr_sel_ram_b4c0_d1 = cbuf_wr_sel_ram_d1[23];
  assign cbuf_p1_wr_sel_ram_b4c1_d1 = cbuf_wr_sel_ram_d1[22];
  assign cbuf_p1_wr_sel_ram_b5c0_d1 = cbuf_wr_sel_ram_d1[21];
  assign cbuf_p1_wr_sel_ram_b5c1_d1 = cbuf_wr_sel_ram_d1[20];
  assign cbuf_p1_wr_sel_ram_b6c0_d1 = cbuf_wr_sel_ram_d1[19];
  assign cbuf_p1_wr_sel_ram_b6c1_d1 = cbuf_wr_sel_ram_d1[18];
  assign cbuf_p1_wr_sel_ram_b7c0_d1 = cbuf_wr_sel_ram_d1[17];
  assign cbuf_p1_wr_sel_ram_b7c1_d1 = cbuf_wr_sel_ram_d1[16];
  assign cbuf_p1_wr_sel_ram_b8c0_d1 = cbuf_wr_sel_ram_d1[15];
  assign cbuf_p1_wr_sel_ram_b8c1_d1 = cbuf_wr_sel_ram_d1[14];
  assign cbuf_p1_wr_sel_ram_b9c0_d1 = cbuf_wr_sel_ram_d1[13];
  assign cbuf_p1_wr_sel_ram_b9c1_d1 = cbuf_wr_sel_ram_d1[12];
  assign cbuf_p2_rd_addr = sc2buf_wmb_rd_addr;
  assign cbuf_p2_rd_c0_data_d4 = cbuf_p2_rd_data_d4[1023:512];
  assign cbuf_p2_rd_c0_data_d6_w = cbuf_p2_rd_c0_data_d5;
  assign cbuf_p2_rd_c0_valid_d5 = cbuf_p2_rd_en_d5;
  assign cbuf_p2_rd_c0_valid_d6_w = cbuf_p2_rd_en_d5;
  assign cbuf_p2_rd_c1_data_d4 = cbuf_p2_rd_data_d4[511:0];
  assign cbuf_p2_rd_c1_data_d6_w = cbuf_p2_rd_c1_data_d5;
  assign cbuf_p2_rd_c1_valid_d5 = cbuf_p2_rd_en_d5;
  assign cbuf_p2_rd_c1_valid_d6_w = cbuf_p2_rd_en_d5;
  assign cbuf_p2_rd_en = sc2buf_wmb_rd_en;
  assign cbuf_p2_rd_en_d3 = cbuf_rd_en_d3[0];
  assign cbuf_p2_rd_en_d4 = cbuf_rd_en_d4[0];
  assign cbuf_p2_rd_sel_ram_b15c0_d3 = cbuf_rd_sel_ram_d3[1];
  assign cbuf_p2_rd_sel_ram_b15c0_w = sc2buf_wmb_rd_en;
  assign cbuf_p2_rd_sel_ram_b15c1_d3 = cbuf_rd_sel_ram_d3[0];
  assign cbuf_p2_rd_sel_ram_b15c1_w = sc2buf_wmb_rd_en;
  assign cbuf_ra_b0c1_w = cbuf_ra_b0c0_w;
  assign cbuf_ra_b10c1_w = cbuf_ra_b10c0_w;
  assign cbuf_ra_b11c1_w = cbuf_ra_b11c0_w;
  assign cbuf_ra_b12c1_w = cbuf_ra_b12c0_w;
  assign cbuf_ra_b13c1_w = cbuf_ra_b13c0_w;
  assign cbuf_ra_b14c1_w = cbuf_ra_b14c0_w;
  assign cbuf_ra_b15c1_w = cbuf_ra_b15c0_w;
  assign cbuf_ra_b1c1_w = cbuf_ra_b1c0_w;
  assign cbuf_ra_b2c1_w = cbuf_ra_b2c0_w;
  assign cbuf_ra_b3c1_w = cbuf_ra_b3c0_w;
  assign cbuf_ra_b4c1_w = cbuf_ra_b4c0_w;
  assign cbuf_ra_b5c1_w = cbuf_ra_b5c0_w;
  assign cbuf_ra_b6c1_w = cbuf_ra_b6c0_w;
  assign cbuf_ra_b7c1_w = cbuf_ra_b7c0_w;
  assign cbuf_ra_b8c1_w = cbuf_ra_b8c0_w;
  assign cbuf_ra_b9c1_w = cbuf_ra_b9c0_w;
  assign cbuf_rd_sel_ram_d1[61] = cbuf_rd_sel_ram_d1[60];
  assign cbuf_rd_sel_ram_d2[61] = cbuf_rd_sel_ram_d2[60];
  assign cbuf_rd_sel_ram_d3[61] = cbuf_rd_sel_ram_d3[60];
  assign cbuf_re_b0c0 = cbuf_re_b0c1;
  assign cbuf_re_b0c0_d2 = cbuf_re_b0c1_d2;
  assign cbuf_re_b0c0_w = cbuf_p0_rd_sel_ram_b0c0_w;
  assign cbuf_re_b0c1_w = cbuf_p0_rd_sel_ram_b0c0_w;
  assign cbuf_re_b10c0 = cbuf_re_b10c1;
  assign cbuf_re_b10c0_d2 = cbuf_re_b10c1_d2;
  assign cbuf_re_b10c1_w = cbuf_re_b10c0_w;
  assign cbuf_re_b11c0 = cbuf_re_b11c1;
  assign cbuf_re_b11c0_d2 = cbuf_re_b11c1_d2;
  assign cbuf_re_b11c1_w = cbuf_re_b11c0_w;
  assign cbuf_re_b12c0 = cbuf_re_b12c1;
  assign cbuf_re_b12c0_d2 = cbuf_re_b12c1_d2;
  assign cbuf_re_b12c1_w = cbuf_re_b12c0_w;
  assign cbuf_re_b13c0 = cbuf_re_b13c1;
  assign cbuf_re_b13c0_d2 = cbuf_re_b13c1_d2;
  assign cbuf_re_b13c1_w = cbuf_re_b13c0_w;
  assign cbuf_re_b14c0 = cbuf_re_b14c1;
  assign cbuf_re_b14c0_d2 = cbuf_re_b14c1_d2;
  assign cbuf_re_b14c1_w = cbuf_re_b14c0_w;
  assign cbuf_re_b15c0 = cbuf_re_b15c1;
  assign cbuf_re_b15c0_d2 = cbuf_re_b15c1_d2;
  assign cbuf_re_b15c1_w = cbuf_re_b15c0_w;
  assign cbuf_re_b1c0 = cbuf_re_b1c1;
  assign cbuf_re_b1c0_d2 = cbuf_re_b1c1_d2;
  assign cbuf_re_b1c1_w = cbuf_re_b1c0_w;
  assign cbuf_re_b2c0 = cbuf_re_b2c1;
  assign cbuf_re_b2c0_d2 = cbuf_re_b2c1_d2;
  assign cbuf_re_b2c1_w = cbuf_re_b2c0_w;
  assign cbuf_re_b3c0 = cbuf_re_b3c1;
  assign cbuf_re_b3c0_d2 = cbuf_re_b3c1_d2;
  assign cbuf_re_b3c1_w = cbuf_re_b3c0_w;
  assign cbuf_re_b4c0 = cbuf_re_b4c1;
  assign cbuf_re_b4c0_d2 = cbuf_re_b4c1_d2;
  assign cbuf_re_b4c1_w = cbuf_re_b4c0_w;
  assign cbuf_re_b5c0 = cbuf_re_b5c1;
  assign cbuf_re_b5c0_d2 = cbuf_re_b5c1_d2;
  assign cbuf_re_b5c1_w = cbuf_re_b5c0_w;
  assign cbuf_re_b6c0 = cbuf_re_b6c1;
  assign cbuf_re_b6c0_d2 = cbuf_re_b6c1_d2;
  assign cbuf_re_b6c1_w = cbuf_re_b6c0_w;
  assign cbuf_re_b7c0 = cbuf_re_b7c1;
  assign cbuf_re_b7c0_d2 = cbuf_re_b7c1_d2;
  assign cbuf_re_b7c1_w = cbuf_re_b7c0_w;
  assign cbuf_re_b8c0 = cbuf_re_b8c1;
  assign cbuf_re_b8c0_d2 = cbuf_re_b8c1_d2;
  assign cbuf_re_b8c1_w = cbuf_re_b8c0_w;
  assign cbuf_re_b9c0 = cbuf_re_b9c1;
  assign cbuf_re_b9c0_d2 = cbuf_re_b9c1_d2;
  assign cbuf_re_b9c1_w = cbuf_re_b9c0_w;
  assign sc2buf_dat_rd_data = cbuf_p0_rd_data_d6;
  assign sc2buf_dat_rd_valid = cbuf_p0_rd_valid_d6;
  assign sc2buf_wmb_rd_data = cbuf_p2_rd_data_d6;
  assign sc2buf_wmb_rd_valid = cbuf_p2_rd_valid_d6;
  assign sc2buf_wt_rd_data = cbuf_p1_rd_data_d6;
  assign sc2buf_wt_rd_valid = cbuf_p1_rd_valid_d6;
endmodule
