module SDP_Y_CORE_chn_mul_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:860" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:861" *)
  output outsig;
  assign outsig = in_0;
endmodule
