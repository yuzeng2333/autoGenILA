module \$paramod\SDP_Y_CVT_mgc_in_wire_v1\rscid=6\width=1 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:78" *)
  output d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:79" *)
  input z;
  assign d = z;
endmodule
