module riscv_core(clk_i, rst_i, mem_d_data_rd_i, mem_d_accept_i, mem_d_ack_i, mem_d_error_i, mem_d_resp_tag_i, mem_i_accept_i, mem_i_valid_i, mem_i_error_i, mem_i_inst_i, intr_i, reset_vector_i, cpu_id_i, mem_d_addr_o, mem_d_data_wr_o, mem_d_rd_o, mem_d_wr_o, mem_d_cacheable_o, mem_d_req_tag_o, mem_d_invalidate_o, mem_d_writeback_o, mem_d_flush_o, mem_i_rd_o, mem_i_flush_o, mem_i_invalidate_o, mem_i_pc_o);
  logic _0000_;
  logic _0001_;
  logic _0002_;
  logic _0003_;
  logic _0004_;
  logic _0005_;
  logic _0006_;
  logic _0007_;
  logic _0008_;
  logic _0009_;
  logic _0010_;
  logic _0011_;
  logic _0012_;
  logic _0013_;
  logic _0014_;
  logic _0015_;
  logic _0016_;
  logic _0017_;
  logic _0018_;
  logic _0019_;
  logic _0020_;
  logic _0021_;
  logic _0022_;
  logic _0023_;
  logic _0024_;
  logic _0025_;
  logic _0026_;
  logic _0027_;
  logic _0028_;
  logic _0029_;
  logic _0030_;
  logic _0031_;
  logic _0032_;
  logic _0033_;
  logic _0034_;
  logic _0035_;
  logic _0036_;
  logic _0037_;
  logic _0038_;
  logic _0039_;
  logic _0040_;
  logic _0041_;
  logic _0042_;
  logic _0043_;
  logic _0044_;
  logic _0045_;
  logic _0046_;
  logic _0047_;
  logic _0048_;
  logic _0049_;
  logic _0050_;
  logic _0051_;
  logic _0052_;
  logic _0053_;
  logic _0054_;
  logic _0055_;
  logic _0056_;
  logic _0057_;
  logic _0058_;
  logic _0059_;
  logic _0060_;
  logic _0061_;
  logic _0062_;
  logic _0063_;
  logic _0064_;
  logic _0065_;
  logic _0066_;
  logic _0067_;
  logic _0068_;
  logic _0069_;
  logic _0070_;
  logic _0071_;
  logic _0072_;
  logic _0073_;
  logic _0074_;
  logic _0075_;
  logic _0076_;
  logic _0077_;
  logic _0078_;
  logic _0079_;
  logic _0080_;
  logic _0081_;
  logic _0082_;
  logic _0083_;
  logic _0084_;
  logic _0085_;
  logic _0086_;
  logic _0087_;
  logic _0088_;
  logic _0089_;
  logic _0090_;
  logic _0091_;
  logic _0092_;
  logic _0093_;
  logic _0094_;
  logic _0095_;
  logic _0096_;
  logic _0097_;
  logic _0098_;
  logic _0099_;
  logic _0100_;
  logic _0101_;
  logic _0102_;
  logic _0103_;
  logic _0104_;
  logic _0105_;
  logic _0106_;
  logic _0107_;
  logic _0108_;
  logic _0109_;
  logic _0110_;
  logic _0111_;
  logic _0112_;
  logic _0113_;
  logic _0114_;
  logic _0115_;
  logic _0116_;
  logic _0117_;
  logic _0118_;
  logic _0119_;
  logic _0120_;
  logic _0121_;
  logic _0122_;
  logic _0123_;
  logic _0124_;
  logic _0125_;
  logic _0126_;
  logic _0127_;
  logic _0128_;
  logic _0129_;
  logic _0130_;
  logic _0131_;
  logic _0132_;
  logic _0133_;
  logic _0134_;
  logic _0135_;
  logic _0136_;
  logic _0137_;
  logic _0138_;
  logic _0139_;
  logic _0140_;
  logic _0141_;
  logic _0142_;
  logic _0143_;
  logic _0144_;
  logic _0145_;
  logic _0146_;
  logic _0147_;
  logic _0148_;
  logic _0149_;
  logic _0150_;
  logic _0151_;
  logic _0152_;
  logic _0153_;
  logic _0154_;
  logic _0155_;
  logic _0156_;
  logic _0157_;
  logic _0158_;
  logic _0159_;
  logic _0160_;
  logic _0161_;
  logic _0162_;
  logic _0163_;
  logic _0164_;
  logic _0165_;
  logic _0166_;
  logic _0167_;
  logic _0168_;
  logic _0169_;
  logic _0170_;
  logic _0171_;
  logic [1:0] _0172_;
  logic [1:0] _0173_;
  logic [1:0] _0174_;
  logic [1:0] _0175_;
  logic [1:0] _0176_;
  logic [1:0] _0177_;
  logic [1:0] _0178_;
  logic [1:0] _0179_;
  logic [1:0] _0180_;
  logic [1:0] _0181_;
  logic _0182_;
  logic _0183_;
  logic _0184_;
  logic _0185_;
  logic _0186_;
  logic _0187_;
  logic _0188_;
  logic _0189_;
  logic _0190_;
  logic _0191_;
  logic [1:0] _0192_;
  logic [1:0] _0193_;
  logic [1:0] _0194_;
  logic [1:0] _0195_;
  logic [1:0] _0196_;
  logic [1:0] _0197_;
  logic [1:0] _0198_;
  logic [1:0] _0199_;
  logic [1:0] _0200_;
  logic [1:0] _0201_;
  logic _0202_;
  logic _0203_;
  logic _0204_;
  logic _0205_;
  logic _0206_;
  logic _0207_;
  logic [31:0] _0208_;
  logic [31:0] _0209_;
  logic [31:0] _0210_;
  logic [31:0] _0211_;
  logic [31:0] _0212_;
  logic [31:0] _0213_;
  logic _0214_;
  logic _0215_;
  logic _0216_;
  logic _0217_;
  logic _0218_;
  logic _0219_;
  logic [63:0] _0220_;
  logic [63:0] _0221_;
  logic [63:0] _0222_;
  logic [63:0] _0223_;
  logic [63:0] _0224_;
  logic [63:0] _0225_;
  logic _0226_;
  logic _0227_;
  logic _0228_;
  logic _0229_;
  logic _0230_;
  logic _0231_;
  logic _0232_;
  logic _0233_;
  logic _0234_;
  logic _0235_;
  logic _0236_;
  logic _0237_;
  logic _0238_;
  logic _0239_;
  logic _0240_;
  logic _0241_;
  logic _0242_;
  logic _0243_;
  logic _0244_;
  logic _0245_;
  logic _0246_;
  logic _0247_;
  logic _0248_;
  logic _0249_;
  logic _0250_;
  logic _0251_;
  logic _0252_;
  logic _0253_;
  logic _0254_;
  logic _0255_;
  logic _0256_;
  logic _0257_;
  logic [1:0] _0258_;
  logic [1:0] _0259_;
  logic [1:0] _0260_;
  logic [1:0] _0261_;
  logic [1:0] _0262_;
  logic [1:0] _0263_;
  logic [1:0] _0264_;
  logic [1:0] _0265_;
  logic [1:0] _0266_;
  logic [1:0] _0267_;
  logic [1:0] _0268_;
  logic [1:0] _0269_;
  logic _0270_;
  logic _0271_;
  logic _0272_;
  logic _0273_;
  logic _0274_;
  logic _0275_;
  logic _0276_;
  logic _0277_;
  logic _0278_;
  logic _0279_;
  logic _0280_;
  logic _0281_;
  logic _0282_;
  logic _0283_;
  logic _0284_;
  logic _0285_;
  logic _0286_;
  logic _0287_;
  logic _0288_;
  logic _0289_;
  logic _0290_;
  logic _0291_;
  logic _0292_;
  logic _0293_;
  logic _0294_;
  logic _0295_;
  logic _0296_;
  logic _0297_;
  logic _0298_;
  logic _0299_;
  logic _0300_;
  logic _0301_;
  logic _0302_;
  logic _0303_;
  logic _0304_;
  logic _0305_;
  logic _0306_;
  logic _0307_;
  logic _0308_;
  logic _0309_;
  logic _0310_;
  logic _0311_;
  logic _0312_;
  logic _0313_;
  logic _0314_;
  logic _0315_;
  logic _0316_;
  logic _0317_;
  logic _0318_;
  logic _0319_;
  logic _0320_;
  logic _0321_;
  logic _0322_;
  logic _0323_;
  logic _0324_;
  logic _0325_;
  logic _0326_;
  logic _0327_;
  logic _0328_;
  logic _0329_;
  logic _0330_;
  logic _0331_;
  logic _0332_;
  logic _0333_;
  logic _0334_;
  logic _0335_;
  logic _0336_;
  logic _0337_;
  logic _0338_;
  logic _0339_;
  logic _0340_;
  logic _0341_;
  logic _0342_;
  logic _0343_;
  logic _0344_;
  logic _0345_;
  logic _0346_;
  logic _0347_;
  logic _0348_;
  logic _0349_;
  logic [1:0] _0350_;
  logic [1:0] _0351_;
  logic [1:0] _0352_;
  logic [1:0] _0353_;
  logic [1:0] _0354_;
  logic [1:0] _0355_;
  logic [1:0] _0356_;
  logic [1:0] _0357_;
  logic [1:0] _0358_;
  logic [1:0] _0359_;
  logic [1:0] _0360_;
  logic [1:0] _0361_;
  logic [1:0] _0362_;
  logic [1:0] _0363_;
  logic [1:0] _0364_;
  logic [1:0] _0365_;
  logic [1:0] _0366_;
  logic [1:0] _0367_;
  logic [1:0] _0368_;
  logic [1:0] _0369_;
  logic [1:0] _0370_;
  logic [1:0] _0371_;
  logic [1:0] _0372_;
  logic [1:0] _0373_;
  logic [1:0] _0374_;
  logic [1:0] _0375_;
  logic [1:0] _0376_;
  logic [1:0] _0377_;
  logic [1:0] _0378_;
  logic [1:0] _0379_;
  logic [1:0] _0380_;
  logic [1:0] _0381_;
  logic [1:0] _0382_;
  logic [1:0] _0383_;
  logic [1:0] _0384_;
  logic [1:0] _0385_;
  logic [1:0] _0386_;
  logic [1:0] _0387_;
  logic [1:0] _0388_;
  logic [1:0] _0389_;
  logic [1:0] _0390_;
  logic [1:0] _0391_;
  logic [1:0] _0392_;
  logic [1:0] _0393_;
  logic [1:0] _0394_;
  logic [1:0] _0395_;
  logic [1:0] _0396_;
  logic [1:0] _0397_;
  logic [1:0] _0398_;
  logic [1:0] _0399_;
  logic [1:0] _0400_;
  logic [1:0] _0401_;
  logic [1:0] _0402_;
  logic [1:0] _0403_;
  logic [1:0] _0404_;
  logic [1:0] _0405_;
  logic [1:0] _0406_;
  logic [1:0] _0407_;
  logic [1:0] _0408_;
  logic [1:0] _0409_;
  logic [1:0] _0410_;
  logic [1:0] _0411_;
  logic [1:0] _0412_;
  logic [1:0] _0413_;
  logic [1:0] _0414_;
  logic [1:0] _0415_;
  logic [1:0] _0416_;
  logic [1:0] _0417_;
  logic [1:0] _0418_;
  logic [1:0] _0419_;
  logic [1:0] _0420_;
  logic [1:0] _0421_;
  logic [1:0] _0422_;
  logic [1:0] _0423_;
  logic [1:0] _0424_;
  logic [1:0] _0425_;
  logic [1:0] _0426_;
  logic [1:0] _0427_;
  logic [1:0] _0428_;
  logic [1:0] _0429_;
  logic _0430_;
  logic _0431_;
  logic _0432_;
  logic _0433_;
  logic _0434_;
  logic _0435_;
  logic _0436_;
  logic _0437_;
  logic _0438_;
  logic _0439_;
  logic _0440_;
  logic _0441_;
  logic _0442_;
  logic _0443_;
  logic _0444_;
  logic _0445_;
  logic _0446_;
  logic _0447_;
  logic _0448_;
  logic _0449_;
  logic _0450_;
  logic _0451_;
  logic _0452_;
  logic _0453_;
  logic _0454_;
  logic _0455_;
  logic _0456_;
  logic _0457_;
  logic _0458_;
  logic _0459_;
  logic _0460_;
  logic _0461_;
  logic _0462_;
  logic _0463_;
  logic _0464_;
  logic _0465_;
  logic _0466_;
  logic _0467_;
  logic _0468_;
  logic _0469_;
  logic _0470_;
  logic _0471_;
  logic _0472_;
  logic _0473_;
  logic _0474_;
  logic _0475_;
  logic _0476_;
  logic _0477_;
  logic _0478_;
  logic _0479_;
  logic _0480_;
  logic _0481_;
  logic _0482_;
  logic _0483_;
  logic _0484_;
  logic _0485_;
  logic _0486_;
  logic _0487_;
  logic _0488_;
  logic _0489_;
  logic _0490_;
  logic _0491_;
  logic _0492_;
  logic _0493_;
  logic _0494_;
  logic _0495_;
  logic _0496_;
  logic _0497_;
  logic _0498_;
  logic _0499_;
  logic _0500_;
  logic _0501_;
  logic _0502_;
  logic _0503_;
  logic _0504_;
  logic _0505_;
  logic _0506_;
  logic _0507_;
  logic _0508_;
  logic _0509_;
  logic _0510_;
  logic _0511_;
  logic _0512_;
  logic _0513_;
  logic _0514_;
  logic _0515_;
  logic _0516_;
  logic _0517_;
  logic _0518_;
  logic _0519_;
  logic _0520_;
  logic _0521_;
  logic _0522_;
  logic _0523_;
  logic _0524_;
  logic _0525_;
  logic _0526_;
  logic _0527_;
  logic _0528_;
  logic _0529_;
  logic _0530_;
  logic _0531_;
  logic _0532_;
  logic _0533_;
  logic _0534_;
  logic _0535_;
  logic _0536_;
  logic _0537_;
  logic _0538_;
  logic _0539_;
  logic _0540_;
  logic _0541_;
  logic _0542_;
  logic _0543_;
  logic _0544_;
  logic _0545_;
  logic _0546_;
  logic _0547_;
  logic _0548_;
  logic _0549_;
  logic _0550_;
  logic _0551_;
  logic _0552_;
  logic _0553_;
  logic _0554_;
  logic _0555_;
  logic _0556_;
  logic _0557_;
  logic _0558_;
  logic _0559_;
  logic _0560_;
  logic _0561_;
  logic _0562_;
  logic _0563_;
  logic _0564_;
  logic _0565_;
  logic _0566_;
  logic _0567_;
  logic _0568_;
  logic _0569_;
  logic _0570_;
  logic _0571_;
  logic _0572_;
  logic _0573_;
  logic _0574_;
  logic _0575_;
  logic _0576_;
  logic _0577_;
  logic _0578_;
  logic _0579_;
  logic _0580_;
  logic _0581_;
  logic _0582_;
  logic _0583_;
  logic _0584_;
  logic _0585_;
  logic _0586_;
  logic _0587_;
  logic _0588_;
  logic _0589_;
  logic _0590_;
  logic _0591_;
  logic _0592_;
  logic _0593_;
  logic _0594_;
  logic _0595_;
  logic _0596_;
  logic _0597_;
  logic _0598_;
  logic _0599_;
  logic _0600_;
  logic _0601_;
  logic _0602_;
  logic _0603_;
  logic _0604_;
  logic _0605_;
  logic _0606_;
  logic _0607_;
  logic _0608_;
  logic _0609_;
  logic _0610_;
  logic _0611_;
  logic _0612_;
  logic _0613_;
  logic _0614_;
  logic _0615_;
  logic _0616_;
  logic _0617_;
  logic _0618_;
  logic _0619_;
  logic _0620_;
  logic _0621_;
  logic _0622_;
  logic _0623_;
  logic _0624_;
  logic _0625_;
  logic _0626_;
  logic _0627_;
  logic _0628_;
  logic _0629_;
  logic _0630_;
  logic _0631_;
  logic _0632_;
  logic _0633_;
  logic _0634_;
  logic _0635_;
  logic _0636_;
  logic _0637_;
  logic _0638_;
  logic _0639_;
  logic _0640_;
  logic _0641_;
  logic _0642_;
  logic _0643_;
  logic _0644_;
  logic _0645_;
  logic _0646_;
  logic _0647_;
  logic _0648_;
  logic _0649_;
  logic _0650_;
  logic _0651_;
  logic _0652_;
  logic _0653_;
  logic _0654_;
  logic _0655_;
  logic _0656_;
  logic _0657_;
  logic _0658_;
  logic _0659_;
  logic _0660_;
  logic _0661_;
  logic _0662_;
  logic _0663_;
  logic _0664_;
  logic _0665_;
  logic _0666_;
  logic _0667_;
  logic _0668_;
  logic _0669_;
  logic _0670_;
  logic _0671_;
  logic _0672_;
  logic _0673_;
  logic _0674_;
  logic _0675_;
  logic _0676_;
  logic _0677_;
  logic _0678_;
  logic _0679_;
  logic _0680_;
  logic _0681_;
  logic _0682_;
  logic _0683_;
  logic _0684_;
  logic _0685_;
  logic _0686_;
  logic _0687_;
  logic _0688_;
  logic _0689_;
  logic _0690_;
  logic _0691_;
  logic _0692_;
  logic _0693_;
  logic _0694_;
  logic _0695_;
  logic _0696_;
  logic _0697_;
  logic _0698_;
  logic _0699_;
  logic _0700_;
  logic _0701_;
  logic _0702_;
  logic _0703_;
  logic _0704_;
  logic _0705_;
  logic _0706_;
  logic _0707_;
  logic _0708_;
  logic _0709_;
  logic _0710_;
  logic _0711_;
  logic _0712_;
  logic _0713_;
  logic _0714_;
  logic _0715_;
  logic _0716_;
  logic _0717_;
  logic _0718_;
  logic _0719_;
  logic _0720_;
  logic _0721_;
  logic _0722_;
  logic _0723_;
  logic _0724_;
  logic _0725_;
  logic _0726_;
  logic _0727_;
  logic _0728_;
  logic _0729_;
  logic _0730_;
  logic _0731_;
  logic _0732_;
  logic _0733_;
  logic _0734_;
  logic _0735_;
  logic _0736_;
  logic _0737_;
  logic _0738_;
  logic _0739_;
  logic _0740_;
  logic _0741_;
  logic _0742_;
  logic _0743_;
  logic _0744_;
  logic _0745_;
  logic _0746_;
  logic _0747_;
  logic _0748_;
  logic _0749_;
  logic _0750_;
  logic _0751_;
  logic _0752_;
  logic _0753_;
  logic _0754_;
  logic _0755_;
  logic _0756_;
  logic _0757_;
  logic _0758_;
  logic _0759_;
  logic _0760_;
  logic _0761_;
  logic _0762_;
  logic _0763_;
  logic _0764_;
  logic _0765_;
  logic _0766_;
  logic _0767_;
  logic _0768_;
  logic _0769_;
  logic _0770_;
  logic _0771_;
  logic _0772_;
  logic _0773_;
  logic _0774_;
  logic _0775_;
  logic _0776_;
  logic _0777_;
  logic _0778_;
  logic _0779_;
  logic _0780_;
  logic _0781_;
  logic _0782_;
  logic _0783_;
  logic _0784_;
  logic _0785_;
  logic _0786_;
  logic _0787_;
  logic _0788_;
  logic _0789_;
  logic _0790_;
  logic _0791_;
  logic _0792_;
  logic _0793_;
  logic _0794_;
  logic _0795_;
  logic _0796_;
  logic _0797_;
  logic _0798_;
  logic _0799_;
  logic _0800_;
  logic _0801_;
  logic _0802_;
  logic _0803_;
  logic _0804_;
  logic _0805_;
  logic _0806_;
  logic _0807_;
  logic _0808_;
  logic _0809_;
  logic _0810_;
  logic _0811_;
  logic _0812_;
  logic _0813_;
  logic _0814_;
  logic _0815_;
  logic _0816_;
  logic _0817_;
  logic _0818_;
  logic _0819_;
  logic _0820_;
  logic _0821_;
  logic _0822_;
  logic _0823_;
  logic _0824_;
  logic _0825_;
  logic _0826_;
  logic _0827_;
  logic _0828_;
  logic _0829_;
  logic _0830_;
  logic _0831_;
  logic _0832_;
  logic _0833_;
  logic _0834_;
  logic _0835_;
  logic _0836_;
  logic _0837_;
  logic _0838_;
  logic _0839_;
  logic _0840_;
  logic _0841_;
  logic _0842_;
  logic _0843_;
  logic _0844_;
  logic _0845_;
  logic _0846_;
  logic _0847_;
  logic _0848_;
  logic _0849_;
  logic _0850_;
  logic _0851_;
  logic _0852_;
  logic _0853_;
  logic _0854_;
  logic _0855_;
  logic _0856_;
  logic _0857_;
  logic _0858_;
  logic _0859_;
  logic _0860_;
  logic _0861_;
  logic _0862_;
  logic _0863_;
  logic _0864_;
  logic _0865_;
  logic _0866_;
  logic _0867_;
  logic _0868_;
  logic _0869_;
  logic _0870_;
  logic _0871_;
  logic _0872_;
  logic _0873_;
  logic _0874_;
  logic _0875_;
  logic _0876_;
  logic _0877_;
  logic _0878_;
  logic _0879_;
  logic _0880_;
  logic _0881_;
  logic _0882_;
  logic _0883_;
  logic _0884_;
  logic _0885_;
  logic _0886_;
  logic _0887_;
  logic _0888_;
  logic _0889_;
  logic _0890_;
  logic _0891_;
  logic _0892_;
  logic _0893_;
  logic _0894_;
  logic _0895_;
  logic _0896_;
  logic _0897_;
  logic _0898_;
  logic _0899_;
  logic _0900_;
  logic _0901_;
  logic _0902_;
  logic _0903_;
  logic _0904_;
  logic _0905_;
  logic _0906_;
  logic _0907_;
  logic _0908_;
  logic _0909_;
  logic _0910_;
  logic _0911_;
  logic _0912_;
  logic _0913_;
  logic _0914_;
  logic _0915_;
  logic _0916_;
  logic _0917_;
  logic _0918_;
  logic _0919_;
  logic _0920_;
  logic _0921_;
  logic _0922_;
  logic _0923_;
  logic _0924_;
  logic _0925_;
  logic _0926_;
  logic _0927_;
  logic _0928_;
  logic _0929_;
  logic _0930_;
  logic _0931_;
  logic _0932_;
  logic _0933_;
  logic _0934_;
  logic _0935_;
  logic _0936_;
  logic _0937_;
  logic _0938_;
  logic _0939_;
  logic _0940_;
  logic _0941_;
  logic _0942_;
  logic _0943_;
  logic _0944_;
  logic _0945_;
  logic _0946_;
  logic _0947_;
  logic _0948_;
  logic _0949_;
  logic _0950_;
  logic _0951_;
  logic _0952_;
  logic _0953_;
  logic _0954_;
  logic _0955_;
  logic _0956_;
  logic _0957_;
  logic _0958_;
  logic _0959_;
  logic _0960_;
  logic _0961_;
  logic _0962_;
  logic _0963_;
  logic _0964_;
  logic _0965_;
  logic _0966_;
  logic _0967_;
  logic _0968_;
  logic _0969_;
  logic _0970_;
  logic _0971_;
  logic _0972_;
  logic _0973_;
  logic _0974_;
  logic _0975_;
  logic _0976_;
  logic _0977_;
  logic _0978_;
  logic _0979_;
  logic _0980_;
  logic _0981_;
  logic _0982_;
  logic _0983_;
  logic _0984_;
  logic _0985_;
  logic _0986_;
  logic _0987_;
  logic _0988_;
  logic _0989_;
  logic _0990_;
  logic _0991_;
  logic _0992_;
  logic _0993_;
  logic _0994_;
  logic _0995_;
  logic _0996_;
  logic _0997_;
  logic _0998_;
  logic _0999_;
  logic _1000_;
  logic _1001_;
  logic _1002_;
  logic _1003_;
  logic _1004_;
  logic _1005_;
  logic _1006_;
  logic _1007_;
  logic _1008_;
  logic _1009_;
  logic _1010_;
  logic _1011_;
  logic _1012_;
  logic _1013_;
  logic _1014_;
  logic _1015_;
  logic _1016_;
  logic _1017_;
  logic _1018_;
  logic _1019_;
  logic _1020_;
  logic _1021_;
  logic _1022_;
  logic _1023_;
  logic _1024_;
  logic _1025_;
  logic _1026_;
  logic _1027_;
  logic _1028_;
  logic _1029_;
  logic _1030_;
  logic _1031_;
  logic _1032_;
  logic _1033_;
  logic _1034_;
  logic _1035_;
  logic _1036_;
  logic _1037_;
  logic _1038_;
  logic _1039_;
  logic _1040_;
  logic _1041_;
  logic _1042_;
  logic _1043_;
  logic _1044_;
  logic _1045_;
  logic _1046_;
  logic _1047_;
  logic _1048_;
  logic _1049_;
  logic _1050_;
  logic _1051_;
  logic _1052_;
  logic _1053_;
  logic [31:0] _1054_;
  logic [31:0] _1055_;
  logic [31:0] _1056_;
  logic [31:0] _1057_;
  logic [31:0] _1058_;
  logic [31:0] _1059_;
  logic [31:0] _1060_;
  logic [31:0] _1061_;
  logic [31:0] _1062_;
  logic [31:0] _1063_;
  logic [31:0] _1064_;
  logic [31:0] _1065_;
  logic [31:0] _1066_;
  logic [31:0] _1067_;
  logic [31:0] _1068_;
  logic [31:0] _1069_;
  logic [31:0] _1070_;
  logic [31:0] _1071_;
  logic [31:0] _1072_;
  logic [31:0] _1073_;
  logic [31:0] _1074_;
  logic [31:0] _1075_;
  logic [31:0] _1076_;
  logic [31:0] _1077_;
  logic [31:0] _1078_;
  logic [31:0] _1079_;
  logic [31:0] _1080_;
  logic [31:0] _1081_;
  logic [31:0] _1082_;
  logic [31:0] _1083_;
  logic [31:0] _1084_;
  logic [31:0] _1085_;
  logic [31:0] _1086_;
  logic [31:0] _1087_;
  logic [31:0] _1088_;
  logic [31:0] _1089_;
  logic [31:0] _1090_;
  logic [31:0] _1091_;
  logic [31:0] _1092_;
  logic [31:0] _1093_;
  logic [31:0] _1094_;
  logic [31:0] _1095_;
  logic [31:0] _1096_;
  logic [31:0] _1097_;
  logic [31:0] _1098_;
  logic [31:0] _1099_;
  logic [31:0] _1100_;
  logic [31:0] _1101_;
  logic _1102_;
  logic _1103_;
  logic _1104_;
  logic _1105_;
  logic _1106_;
  logic _1107_;
  logic _1108_;
  logic _1109_;
  logic _1110_;
  logic _1111_;
  logic _1112_;
  logic _1113_;
  logic _1114_;
  logic _1115_;
  logic _1116_;
  logic _1117_;
  logic _1118_;
  logic _1119_;
  logic _1120_;
  logic _1121_;
  logic _1122_;
  logic _1123_;
  logic _1124_;
  logic _1125_;
  logic _1126_;
  logic _1127_;
  logic _1128_;
  logic _1129_;
  logic _1130_;
  logic _1131_;
  logic _1132_;
  logic _1133_;
  logic _1134_;
  logic _1135_;
  logic _1136_;
  logic _1137_;
  logic _1138_;
  logic _1139_;
  logic _1140_;
  logic _1141_;
  logic _1142_;
  logic _1143_;
  logic _1144_;
  logic _1145_;
  logic _1146_;
  logic _1147_;
  logic _1148_;
  logic _1149_;
  logic _1150_;
  logic _1151_;
  logic _1152_;
  logic _1153_;
  logic _1154_;
  logic _1155_;
  logic _1156_;
  logic _1157_;
  logic _1158_;
  logic _1159_;
  logic _1160_;
  logic _1161_;
  logic _1162_;
  logic _1163_;
  logic _1164_;
  logic _1165_;
  logic _1166_;
  logic _1167_;
  logic _1168_;
  logic _1169_;
  logic _1170_;
  logic _1171_;
  logic _1172_;
  logic _1173_;
  logic _1174_;
  logic _1175_;
  logic _1176_;
  logic _1177_;
  logic _1178_;
  logic _1179_;
  logic _1180_;
  logic _1181_;
  logic [31:0] _1182_;
  logic [31:0] _1183_;
  logic [31:0] _1184_;
  logic [31:0] _1185_;
  logic [31:0] _1186_;
  logic [31:0] _1187_;
  logic [31:0] _1188_;
  logic [31:0] _1189_;
  logic [31:0] _1190_;
  logic [31:0] _1191_;
  logic [31:0] _1192_;
  logic [31:0] _1193_;
  logic [31:0] _1194_;
  logic [31:0] _1195_;
  logic [31:0] _1196_;
  logic [31:0] _1197_;
  logic [31:0] _1198_;
  logic [31:0] _1199_;
  logic [31:0] _1200_;
  logic [31:0] _1201_;
  logic [31:0] _1202_;
  logic [31:0] _1203_;
  logic [31:0] _1204_;
  logic [31:0] _1205_;
  logic [31:0] _1206_;
  logic [31:0] _1207_;
  logic [31:0] _1208_;
  logic [31:0] _1209_;
  logic [31:0] _1210_;
  logic [31:0] _1211_;
  logic [31:0] _1212_;
  logic [31:0] _1213_;
  logic [31:0] _1214_;
  logic [31:0] _1215_;
  logic [31:0] _1216_;
  logic [31:0] _1217_;
  logic [31:0] _1218_;
  logic [31:0] _1219_;
  logic [31:0] _1220_;
  logic [31:0] _1221_;
  logic [31:0] _1222_;
  logic [31:0] _1223_;
  logic [31:0] _1224_;
  logic [31:0] _1225_;
  logic [31:0] _1226_;
  logic [31:0] _1227_;
  logic [31:0] _1228_;
  logic [31:0] _1229_;
  logic [31:0] _1230_;
  logic [31:0] _1231_;
  logic [31:0] _1232_;
  logic [31:0] _1233_;
  logic [31:0] _1234_;
  logic [31:0] _1235_;
  logic [31:0] _1236_;
  logic [31:0] _1237_;
  logic [31:0] _1238_;
  logic [31:0] _1239_;
  logic [31:0] _1240_;
  logic [31:0] _1241_;
  logic [31:0] _1242_;
  logic [31:0] _1243_;
  logic [31:0] _1244_;
  logic [31:0] _1245_;
  logic [31:0] _1246_;
  logic [31:0] _1247_;
  logic [31:0] _1248_;
  logic [31:0] _1249_;
  logic [31:0] _1250_;
  logic [31:0] _1251_;
  logic [31:0] _1252_;
  logic [31:0] _1253_;
  logic [31:0] _1254_;
  logic [31:0] _1255_;
  logic [31:0] _1256_;
  logic [31:0] _1257_;
  logic [31:0] _1258_;
  logic [31:0] _1259_;
  logic [31:0] _1260_;
  logic [31:0] _1261_;
  logic [31:0] _1262_;
  logic [31:0] _1263_;
  logic [31:0] _1264_;
  logic [31:0] _1265_;
  logic [31:0] _1266_;
  logic [31:0] _1267_;
  logic [31:0] _1268_;
  logic [31:0] _1269_;
  logic [31:0] _1270_;
  logic [31:0] _1271_;
  logic [31:0] _1272_;
  logic [31:0] _1273_;
  logic [31:0] _1274_;
  logic [31:0] _1275_;
  logic [31:0] _1276_;
  logic [31:0] _1277_;
  logic [31:0] _1278_;
  logic [31:0] _1279_;
  logic [31:0] _1280_;
  logic [31:0] _1281_;
  logic [31:0] _1282_;
  logic [31:0] _1283_;
  logic [31:0] _1284_;
  logic [31:0] _1285_;
  logic [31:0] _1286_;
  logic [31:0] _1287_;
  logic [31:0] _1288_;
  logic [31:0] _1289_;
  logic [31:0] _1290_;
  logic [31:0] _1291_;
  logic [31:0] _1292_;
  logic [31:0] _1293_;
  logic [31:0] _1294_;
  logic [31:0] _1295_;
  logic [31:0] _1296_;
  logic [31:0] _1297_;
  logic [31:0] _1298_;
  logic [31:0] _1299_;
  logic [31:0] _1300_;
  logic [31:0] _1301_;
  logic [31:0] _1302_;
  logic [31:0] _1303_;
  logic [31:0] _1304_;
  logic [31:0] _1305_;
  logic [31:0] _1306_;
  logic [31:0] _1307_;
  logic [31:0] _1308_;
  logic [31:0] _1309_;
  logic _1310_;
  logic _1311_;
  logic _1312_;
  logic _1313_;
  logic _1314_;
  logic _1315_;
  logic _1316_;
  logic _1317_;
  logic _1318_;
  logic _1319_;
  logic _1320_;
  logic _1321_;
  logic _1322_;
  logic _1323_;
  logic _1324_;
  logic _1325_;
  logic _1326_;
  logic _1327_;
  logic _1328_;
  logic _1329_;
  logic _1330_;
  logic _1331_;
  logic _1332_;
  logic _1333_;
  logic _1334_;
  logic _1335_;
  logic _1336_;
  logic _1337_;
  logic _1338_;
  logic _1339_;
  logic _1340_;
  logic _1341_;
  logic _1342_;
  logic _1343_;
  logic _1344_;
  logic _1345_;
  logic _1346_;
  logic _1347_;
  logic _1348_;
  logic _1349_;
  logic _1350_;
  logic _1351_;
  logic _1352_;
  logic _1353_;
  logic _1354_;
  logic _1355_;
  logic _1356_;
  logic _1357_;
  logic _1358_;
  logic _1359_;
  logic _1360_;
  logic _1361_;
  logic _1362_;
  logic _1363_;
  logic _1364_;
  logic _1365_;
  logic _1366_;
  logic _1367_;
  logic _1368_;
  logic _1369_;
  logic _1370_;
  logic _1371_;
  logic _1372_;
  logic _1373_;
  logic _1374_;
  logic _1375_;
  logic _1376_;
  logic _1377_;
  logic _1378_;
  logic _1379_;
  logic _1380_;
  logic _1381_;
  logic _1382_;
  logic _1383_;
  logic _1384_;
  logic _1385_;
  logic _1386_;
  logic _1387_;
  logic _1388_;
  logic _1389_;
  logic [31:0] _1390_;
  logic [31:0] _1391_;
  logic [31:0] _1392_;
  logic [31:0] _1393_;
  logic [31:0] _1394_;
  logic [31:0] _1395_;
  logic [31:0] _1396_;
  logic [31:0] _1397_;
  logic [31:0] _1398_;
  logic [31:0] _1399_;
  logic [31:0] _1400_;
  logic [31:0] _1401_;
  logic [31:0] _1402_;
  logic [31:0] _1403_;
  logic [31:0] _1404_;
  logic [31:0] _1405_;
  logic [31:0] _1406_;
  logic [31:0] _1407_;
  logic [31:0] _1408_;
  logic [31:0] _1409_;
  logic [31:0] _1410_;
  logic [31:0] _1411_;
  logic [31:0] _1412_;
  logic [31:0] _1413_;
  logic [31:0] _1414_;
  logic [31:0] _1415_;
  logic [31:0] _1416_;
  logic [31:0] _1417_;
  logic [31:0] _1418_;
  logic [31:0] _1419_;
  logic [31:0] _1420_;
  logic [31:0] _1421_;
  logic [31:0] _1422_;
  logic [31:0] _1423_;
  logic [31:0] _1424_;
  logic [31:0] _1425_;
  logic [31:0] _1426_;
  logic [31:0] _1427_;
  logic [31:0] _1428_;
  logic [31:0] _1429_;
  logic [31:0] _1430_;
  logic [31:0] _1431_;
  logic [31:0] _1432_;
  logic [31:0] _1433_;
  logic [31:0] _1434_;
  logic [31:0] _1435_;
  logic [31:0] _1436_;
  logic [31:0] _1437_;
  logic [31:0] _1438_;
  logic [31:0] _1439_;
  logic [31:0] _1440_;
  logic [31:0] _1441_;
  logic [31:0] _1442_;
  logic [31:0] _1443_;
  logic [31:0] _1444_;
  logic [31:0] _1445_;
  logic [31:0] _1446_;
  logic [31:0] _1447_;
  logic [31:0] _1448_;
  logic [31:0] _1449_;
  logic [31:0] _1450_;
  logic [31:0] _1451_;
  logic [31:0] _1452_;
  logic [31:0] _1453_;
  logic [31:0] _1454_;
  logic [31:0] _1455_;
  logic [31:0] _1456_;
  logic [31:0] _1457_;
  logic [31:0] _1458_;
  logic [31:0] _1459_;
  logic [31:0] _1460_;
  logic [31:0] _1461_;
  logic [31:0] _1462_;
  logic [31:0] _1463_;
  logic [31:0] _1464_;
  logic [31:0] _1465_;
  logic [31:0] _1466_;
  logic [31:0] _1467_;
  logic [31:0] _1468_;
  logic [31:0] _1469_;
  logic [31:0] _1470_;
  logic [31:0] _1471_;
  logic [31:0] _1472_;
  logic [31:0] _1473_;
  logic [31:0] _1474_;
  logic [31:0] _1475_;
  logic _1476_;
  logic _1477_;
  logic _1478_;
  logic _1479_;
  logic _1480_;
  logic _1481_;
  logic _1482_;
  logic _1483_;
  logic _1484_;
  logic _1485_;
  logic _1486_;
  logic _1487_;
  logic _1488_;
  logic _1489_;
  logic _1490_;
  logic _1491_;
  logic _1492_;
  logic _1493_;
  logic _1494_;
  logic _1495_;
  logic _1496_;
  logic _1497_;
  logic _1498_;
  logic _1499_;
  logic _1500_;
  logic _1501_;
  logic _1502_;
  logic _1503_;
  logic _1504_;
  logic _1505_;
  logic _1506_;
  logic _1507_;
  logic _1508_;
  logic _1509_;
  logic _1510_;
  logic _1511_;
  logic _1512_;
  logic _1513_;
  logic _1514_;
  logic _1515_;
  logic _1516_;
  logic _1517_;
  logic _1518_;
  logic _1519_;
  logic _1520_;
  logic _1521_;
  logic _1522_;
  logic _1523_;
  logic _1524_;
  logic _1525_;
  logic _1526_;
  logic _1527_;
  logic _1528_;
  logic _1529_;
  logic _1530_;
  logic _1531_;
  logic _1532_;
  logic _1533_;
  logic _1534_;
  logic _1535_;
  logic _1536_;
  logic _1537_;
  logic _1538_;
  logic _1539_;
  logic _1540_;
  logic _1541_;
  logic _1542_;
  logic _1543_;
  logic _1544_;
  logic _1545_;
  logic _1546_;
  logic _1547_;
  logic _1548_;
  logic _1549_;
  logic _1550_;
  logic _1551_;
  logic _1552_;
  logic _1553_;
  logic _1554_;
  logic _1555_;
  logic [31:0] _1556_;
  logic [31:0] _1557_;
  logic [31:0] _1558_;
  logic [31:0] _1559_;
  logic [31:0] _1560_;
  logic [31:0] _1561_;
  logic [31:0] _1562_;
  logic [31:0] _1563_;
  logic [31:0] _1564_;
  logic [31:0] _1565_;
  logic [31:0] _1566_;
  logic [31:0] _1567_;
  logic [31:0] _1568_;
  logic [31:0] _1569_;
  logic [31:0] _1570_;
  logic [31:0] _1571_;
  logic [31:0] _1572_;
  logic [31:0] _1573_;
  logic [31:0] _1574_;
  logic [31:0] _1575_;
  logic [31:0] _1576_;
  logic [31:0] _1577_;
  logic [31:0] _1578_;
  logic [31:0] _1579_;
  logic [31:0] _1580_;
  logic [31:0] _1581_;
  logic [31:0] _1582_;
  logic [31:0] _1583_;
  logic [31:0] _1584_;
  logic [31:0] _1585_;
  logic [31:0] _1586_;
  logic [31:0] _1587_;
  logic [31:0] _1588_;
  logic [31:0] _1589_;
  logic [31:0] _1590_;
  logic [31:0] _1591_;
  logic [31:0] _1592_;
  logic [31:0] _1593_;
  logic [31:0] _1594_;
  logic [31:0] _1595_;
  logic [31:0] _1596_;
  logic [31:0] _1597_;
  logic [31:0] _1598_;
  logic [31:0] _1599_;
  logic [31:0] _1600_;
  logic [31:0] _1601_;
  logic [31:0] _1602_;
  logic [31:0] _1603_;
  logic [31:0] _1604_;
  logic [31:0] _1605_;
  logic [31:0] _1606_;
  logic [31:0] _1607_;
  logic [31:0] _1608_;
  logic [31:0] _1609_;
  logic [31:0] _1610_;
  logic [31:0] _1611_;
  logic [31:0] _1612_;
  logic [31:0] _1613_;
  logic [31:0] _1614_;
  logic [31:0] _1615_;
  logic [31:0] _1616_;
  logic [31:0] _1617_;
  logic [31:0] _1618_;
  logic [31:0] _1619_;
  logic [31:0] _1620_;
  logic [31:0] _1621_;
  logic [31:0] _1622_;
  logic [31:0] _1623_;
  logic [31:0] _1624_;
  logic [31:0] _1625_;
  logic [31:0] _1626_;
  logic [31:0] _1627_;
  logic [31:0] _1628_;
  logic [31:0] _1629_;
  logic [31:0] _1630_;
  logic [31:0] _1631_;
  logic [31:0] _1632_;
  logic [31:0] _1633_;
  logic [31:0] _1634_;
  logic [31:0] _1635_;
  logic _1636_;
  logic _1637_;
  logic _1638_;
  logic _1639_;
  logic _1640_;
  logic _1641_;
  logic [35:0] _1642_;
  logic [35:0] _1643_;
  logic [35:0] _1644_;
  logic [35:0] _1645_;
  logic [35:0] _1646_;
  logic [35:0] _1647_;
  logic _1648_;
  logic [31:0] _1649_;
  logic [31:0] _1650_;
  logic [5:0] _1651_;
  logic _1652_;
  logic [31:0] _1653_;
  logic _1654_;
  logic _1655_;
  logic _1656_;
  logic [5:0] _1657_;
  logic [31:0] _1658_;
  logic [31:0] _1659_;
  logic [31:0] _1660_;
  logic [31:0] _1661_;
  logic _1662_;
  logic [31:0] _1663_;
  logic _1664_;
  logic _1665_;
  logic _1666_;
  logic _1667_;
  logic _1668_;
  logic _1669_;
  logic _1670_;
  logic _1671_;
  logic _1672_;
  logic _1673_;
  logic _1674_;
  logic _1675_;
  logic _1676_;
  logic _1677_;
  logic _1678_;
  logic _1679_;
  logic _1680_;
  logic _1681_;
  logic _1682_;
  logic [31:0] _1683_;
  logic _1684_;
  logic _1685_;
  logic _1686_;
  logic _1687_;
  logic _1688_;
  logic _1689_;
  logic _1690_;
  logic _1691_;
  logic [31:0] _1692_;
  logic [31:0] _1693_;
  logic _1694_;
  logic [5:0] _1695_;
  logic [5:0] _1696_;
  logic [5:0] _1697_;
  logic [5:0] _1698_;
  logic [5:0] _1699_;
  logic [5:0] _1700_;
  logic [31:0] _1701_;
  logic [31:0] _1702_;
  logic [31:0] _1703_;
  logic [31:0] _1704_;
  logic [31:0] _1705_;
  logic [31:0] _1706_;
  logic _1707_;
  logic _1708_;
  logic [31:0] _1709_;
  logic [31:0] _1710_;
  logic [31:0] _1711_;
  logic [31:0] _1712_;
  logic [31:0] _1713_;
  logic [31:0] _1714_;
  logic _1715_;
  logic [31:0] _1716_;
  logic [31:0] _1717_;
  logic [31:0] _1718_;
  logic [31:0] _1719_;
  logic [1:0] _1720_;
  logic _1721_;
  logic [1:0] _1722_;
  logic [1:0] _1723_;
  logic [31:0] _1724_;
  logic [31:0] _1725_;
  logic [31:0] _1726_;
  logic _1727_;
  logic [31:0] _1728_;
  logic [31:0] _1729_;
  logic [31:0] _1730_;
  logic [31:0] _1731_;
  logic [31:0] _1732_;
  logic [31:0] _1733_;
  logic [31:0] _1734_;
  logic [31:0] _1735_;
  logic _1736_;
  logic [31:0] _1737_;
  logic [31:0] _1738_;
  logic [31:0] _1739_;
  logic [31:0] _1740_;
  logic _1741_;
  logic [31:0] _1742_;
  logic [31:0] _1743_;
  logic [31:0] _1744_;
  logic [31:0] _1745_;
  logic _1746_;
  logic _1747_;
  logic [31:0] _1748_;
  logic [31:0] _1749_;
  logic [31:0] _1750_;
  logic _1751_;
  logic [31:0] _1752_;
  logic _1753_;
  logic [31:0] _1754_;
  logic [31:0] _1755_;
  logic [31:0] _1756_;
  logic [31:0] _1757_;
  logic [31:0] _1758_;
  logic [1:0] _1759_;
  logic _1760_;
  logic [31:0] _1761_;
  logic [31:0] _1762_;
  logic [31:0] _1763_;
  logic [31:0] _1764_;
  logic [1:0] _1765_;
  logic [31:0] _1766_;
  logic _1767_;
  logic [31:0] _1768_;
  logic [31:0] _1769_;
  logic _1770_;
  logic _1771_;
  logic [31:0] _1772_;
  logic _1773_;
  logic [31:0] _1774_;
  logic [31:0] _1775_;
  logic [31:0] _1776_;
  logic [31:0] _1777_;
  logic [31:0] _1778_;
  logic [31:0] _1779_;
  logic [31:0] _1780_;
  logic [31:0] _1781_;
  logic [31:0] _1782_;
  logic [5:0] _1783_;
  logic [31:0] _1784_;
  logic [31:0] _1785_;
  logic [31:0] _1786_;
  logic [31:0] _1787_;
  logic [31:0] _1788_;
  logic [31:0] _1789_;
  logic [31:0] _1790_;
  logic [31:0] _1791_;
  logic _1792_;
  logic _1793_;
  logic _1794_;
  logic _1795_;
  logic _1796_;
  logic _1797_;
  logic _1798_;
  logic _1799_;
  logic _1800_;
  logic _1801_;
  logic _1802_;
  logic _1803_;
  logic _1804_;
  logic _1805_;
  logic _1806_;
  logic _1807_;
  logic _1808_;
  logic _1809_;
  logic _1810_;
  logic _1811_;
  logic _1812_;
  logic _1813_;
  logic _1814_;
  logic _1815_;
  logic _1816_;
  logic [31:0] _1817_;
  logic [31:0] _1818_;
  logic [31:0] _1819_;
  logic _1820_;
  logic _1821_;
  logic _1822_;
  logic _1823_;
  logic _1824_;
  logic _1825_;
  logic _1826_;
  logic _1827_;
  logic _1828_;
  logic [6:0] _1829_;
  logic _1830_;
  logic [2:0] _1831_;
  logic _1832_;
  logic _1833_;
  logic _1834_;
  logic [1:0] _1835_;
  logic _1836_;
  logic _1837_;
  logic _1838_;
  logic _1839_;
  logic _1840_;
  logic _1841_;
  logic _1842_;
  logic _1843_;
  logic _1844_;
  logic _1845_;
  logic [1:0] _1846_;
  logic _1847_;
  logic _1848_;
  logic [31:0] _1849_;
  logic [31:0] _1850_;
  logic _1851_;
  logic _1852_;
  logic [31:0] _1853_;
  logic [62:0] _1854_;
  logic _1855_;
  logic [31:0] _1856_;
  logic [31:0] _1857_;
  logic _1858_;
  logic _1859_;
  logic _1860_;
  logic _1861_;
  logic [31:0] _1862_;
  logic [31:0] _1863_;
  logic _1864_;
  logic [31:0] _1865_;
  logic [31:0] _1866_;
  logic _1867_;
  logic _1868_;
  logic _1869_;
  logic _1870_;
  logic _1871_;
  logic _1872_;
  logic _1873_;
  logic _1874_;
  logic _1875_;
  logic _1876_;
  logic _1877_;
  logic _1878_;
  logic _1879_;
  logic _1880_;
  logic _1881_;
  logic _1882_;
  logic _1883_;
  logic _1884_;
  logic _1885_;
  logic _1886_;
  logic _1887_;
  logic [31:0] _1888_;
  logic [31:0] _1889_;
  logic [31:0] _1890_;
  logic [31:0] _1891_;
  logic [31:0] _1892_;
  logic [31:0] _1893_;
  logic _1894_;
  logic _1895_;
  logic _1896_;
  logic _1897_;
  logic _1898_;
  logic _1899_;
  logic _1900_;
  logic _1901_;
  logic [31:0] _1902_;
  logic [31:0] _1903_;
  logic [31:0] _1904_;
  logic [31:0] _1905_;
  logic _1906_;
  logic _1907_;
  logic _1908_;
  logic _1909_;
  logic _1910_;
  logic _1911_;
  logic [31:0] _1912_;
  logic [31:0] _1913_;
  logic [31:0] _1914_;
  logic [31:0] _1915_;
  logic [31:0] _1916_;
  logic [31:0] _1917_;
  logic [31:0] _1918_;
  logic [31:0] _1919_;
  logic [31:0] _1920_;
  logic [62:0] _1921_;
  logic [62:0] _1922_;
  logic [62:0] _1923_;
  logic [62:0] _1924_;
  logic [62:0] _1925_;
  logic [31:0] _1926_;
  logic [31:0] _1927_;
  logic [31:0] _1928_;
  logic [31:0] _1929_;
  logic [31:0] _1930_;
  logic [31:0] _1931_;
  logic _1932_;
  logic _1933_;
  logic [31:0] _1934_;
  logic [31:0] _1935_;
  logic [31:0] _1936_;
  logic _1937_;
  logic _1938_;
  logic _1939_;
  logic _1940_;
  logic _1941_;
  logic [31:0] _1942_;
  logic [31:0] _1943_;
  logic [31:0] _1944_;
  logic [3:0] _1945_;
  logic [31:0] _1946_;
  logic [31:0] _1947_;
  logic [3:0] _1948_;
  logic [31:0] _1949_;
  logic [31:0] _1950_;
  logic [3:0] _1951_;
  logic [31:0] _1952_;
  logic [31:0] _1953_;
  logic [3:0] _1954_;
  logic [31:0] _1955_;
  logic [31:0] _1956_;
  logic [3:0] _1957_;
  logic [31:0] _1958_;
  logic [31:0] _1959_;
  logic [3:0] _1960_;
  logic [31:0] _1961_;
  logic [31:0] _1962_;
  logic [3:0] _1963_;
  logic [31:0] _1964_;
  logic [31:0] _1965_;
  logic [3:0] _1966_;
  logic [31:0] _1967_;
  logic [31:0] _1968_;
  logic [3:0] _1969_;
  logic [31:0] _1970_;
  logic [31:0] _1971_;
  logic [3:0] _1972_;
  logic [31:0] _1973_;
  logic [31:0] _1974_;
  logic [3:0] _1975_;
  logic [31:0] _1976_;
  logic [31:0] _1977_;
  logic [3:0] _1978_;
  logic [31:0] _1979_;
  logic [31:0] _1980_;
  logic [2:0] _1981_;
  logic [31:0] _1982_;
  logic [3:0] _1983_;
  logic [31:0] _1984_;
  logic [31:0] _1985_;
  logic _1986_;
  logic _1987_;
  logic _1988_;
  logic _1989_;
  logic _1990_;
  logic [31:0] _1991_;
  logic [3:0] _1992_;
  logic [31:0] _1993_;
  logic [31:0] _1994_;
  logic _1995_;
  logic _1996_;
  logic [3:0] _1997_;
  logic [31:0] _1998_;
  logic [31:0] _1999_;
  logic _2000_;
  logic _2001_;
  logic [3:0] _2002_;
  logic [31:0] _2003_;
  logic [31:0] _2004_;
  logic _2005_;
  logic _2006_;
  logic _2007_;
  logic [3:0] _2008_;
  logic [31:0] _2009_;
  logic [31:0] _2010_;
  logic _2011_;
  logic _2012_;
  logic _2013_;
  logic [3:0] _2014_;
  logic [31:0] _2015_;
  logic [31:0] _2016_;
  logic _2017_;
  logic _2018_;
  logic [3:0] _2019_;
  logic [31:0] _2020_;
  logic [31:0] _2021_;
  logic _2022_;
  logic _2023_;
  logic [3:0] _2024_;
  logic [31:0] _2025_;
  logic [31:0] _2026_;
  logic [31:0] _2027_;
  logic [31:0] _2028_;
  logic [31:0] _2029_;
  logic [31:0] _2030_;
  logic [31:0] _2031_;
  logic [31:0] _2032_;
  logic [31:0] _2033_;
  logic [31:0] _2034_;
  logic _2035_;
  logic _2036_;
  logic _2037_;
  logic _2038_;
  logic _2039_;
  logic _2040_;
  logic _2041_;
  logic _2042_;
  logic _2043_;
  logic _2044_;
  logic _2045_;
  logic _2046_;
  logic _2047_;
  logic _2048_;
  logic _2049_;
  logic _2050_;
  logic _2051_;
  logic _2052_;
  logic _2053_;
  logic _2054_;
  logic _2055_;
  logic _2056_;
  logic _2057_;
  logic _2058_;
  logic _2059_;
  logic _2060_;
  logic _2061_;
  logic _2062_;
  logic _2063_;
  logic _2064_;
  logic _2065_;
  logic _2066_;
  logic _2067_;
  logic _2068_;
  logic _2069_;
  logic _2070_;
  logic _2071_;
  logic _2072_;
  logic _2073_;
  logic _2074_;
  logic _2075_;
  logic _2076_;
  logic _2077_;
  logic _2078_;
  logic _2079_;
  logic _2080_;
  logic _2081_;
  logic _2082_;
  logic _2083_;
  logic _2084_;
  logic _2085_;
  logic _2086_;
  logic _2087_;
  logic _2088_;
  logic _2089_;
  logic _2090_;
  logic [31:0] _2091_;
  logic [31:0] _2092_;
  logic _2093_;
  logic _2094_;
  logic [31:0] _2095_;
  logic [31:0] _2096_;
  logic [31:0] _2097_;
  logic [31:0] _2098_;
  logic [31:0] _2099_;
  logic [31:0] _2100_;
  logic [31:0] _2101_;
  logic [31:0] _2102_;
  logic [31:0] _2103_;
  logic [31:0] _2104_;
  logic [31:0] _2105_;
  logic [31:0] _2106_;
  logic [31:0] _2107_;
  logic [15:0] _2108_;
  logic [31:0] _2109_;
  logic _2110_;
  logic [31:0] _2111_;
  logic [31:0] _2112_;
  logic [1:0] _2113_;
  logic [31:0] _2114_;
  logic _2115_;
  logic _2116_;
  logic _2117_;
  logic _2118_;
  logic [31:0] _2119_;
  logic _2120_;
  logic _2121_;
  logic _2122_;
  logic _2123_;
  logic _2124_;
  logic _2125_;
  logic _2126_;
  logic _2127_;
  logic _2128_;
  logic [31:0] _2129_;
  logic [31:0] _2130_;
  logic [31:0] _2131_;
  logic _2132_;
  logic _2133_;
  logic _2134_;
  logic _2135_;
  logic _2136_;
  logic [31:0] _2137_;
  logic [31:0] _2138_;
  logic [31:0] _2139_;
  logic [3:0] _2140_;
  logic [31:0] _2141_;
  logic [31:0] _2142_;
  logic [3:0] _2143_;
  logic [31:0] _2144_;
  logic [31:0] _2145_;
  logic [3:0] _2146_;
  logic [31:0] _2147_;
  logic [31:0] _2148_;
  logic [3:0] _2149_;
  logic [31:0] _2150_;
  logic [31:0] _2151_;
  logic [3:0] _2152_;
  logic [31:0] _2153_;
  logic [31:0] _2154_;
  logic [3:0] _2155_;
  logic [31:0] _2156_;
  logic [31:0] _2157_;
  logic [3:0] _2158_;
  logic [31:0] _2159_;
  logic [31:0] _2160_;
  logic [3:0] _2161_;
  logic [31:0] _2162_;
  logic [31:0] _2163_;
  logic [3:0] _2164_;
  logic [31:0] _2165_;
  logic [31:0] _2166_;
  logic [3:0] _2167_;
  logic [31:0] _2168_;
  logic [31:0] _2169_;
  logic [3:0] _2170_;
  logic [31:0] _2171_;
  logic [31:0] _2172_;
  logic [3:0] _2173_;
  logic [31:0] _2174_;
  logic [31:0] _2175_;
  logic [2:0] _2176_;
  logic [31:0] _2177_;
  logic [3:0] _2178_;
  logic [31:0] _2179_;
  logic [31:0] _2180_;
  logic _2181_;
  logic _2182_;
  logic _2183_;
  logic _2184_;
  logic _2185_;
  logic [31:0] _2186_;
  logic [3:0] _2187_;
  logic [31:0] _2188_;
  logic [31:0] _2189_;
  logic _2190_;
  logic _2191_;
  logic [3:0] _2192_;
  logic [31:0] _2193_;
  logic [31:0] _2194_;
  logic _2195_;
  logic _2196_;
  logic [3:0] _2197_;
  logic [31:0] _2198_;
  logic [31:0] _2199_;
  logic _2200_;
  logic _2201_;
  logic _2202_;
  logic [3:0] _2203_;
  logic [31:0] _2204_;
  logic [31:0] _2205_;
  logic _2206_;
  logic _2207_;
  logic _2208_;
  logic [3:0] _2209_;
  logic [31:0] _2210_;
  logic [31:0] _2211_;
  logic _2212_;
  logic _2213_;
  logic [3:0] _2214_;
  logic [31:0] _2215_;
  logic [31:0] _2216_;
  logic _2217_;
  logic _2218_;
  logic [3:0] _2219_;
  logic [31:0] _2220_;
  logic [31:0] _2221_;
  logic [31:0] _2222_;
  logic [31:0] _2223_;
  logic [31:0] _2224_;
  logic [31:0] _2225_;
  logic [31:0] _2226_;
  logic [31:0] _2227_;
  logic [31:0] _2228_;
  logic [31:0] _2229_;
  logic _2230_;
  logic _2231_;
  logic _2232_;
  logic _2233_;
  logic _2234_;
  logic _2235_;
  logic _2236_;
  logic _2237_;
  logic _2238_;
  logic _2239_;
  logic _2240_;
  logic _2241_;
  logic _2242_;
  logic _2243_;
  logic _2244_;
  logic _2245_;
  logic _2246_;
  logic _2247_;
  logic _2248_;
  logic _2249_;
  logic _2250_;
  logic _2251_;
  logic _2252_;
  logic _2253_;
  logic _2254_;
  logic _2255_;
  logic _2256_;
  logic _2257_;
  logic _2258_;
  logic _2259_;
  logic _2260_;
  logic _2261_;
  logic _2262_;
  logic _2263_;
  logic _2264_;
  logic _2265_;
  logic _2266_;
  logic _2267_;
  logic _2268_;
  logic _2269_;
  logic _2270_;
  logic _2271_;
  logic _2272_;
  logic _2273_;
  logic _2274_;
  logic _2275_;
  logic _2276_;
  logic _2277_;
  logic _2278_;
  logic _2279_;
  logic _2280_;
  logic _2281_;
  logic _2282_;
  logic _2283_;
  logic _2284_;
  logic _2285_;
  logic [31:0] _2286_;
  logic [31:0] _2287_;
  logic _2288_;
  logic _2289_;
  logic [31:0] _2290_;
  logic [31:0] _2291_;
  logic [31:0] _2292_;
  logic [31:0] _2293_;
  logic [31:0] _2294_;
  logic [31:0] _2295_;
  logic [31:0] _2296_;
  logic [31:0] _2297_;
  logic [31:0] _2298_;
  logic [31:0] _2299_;
  logic [31:0] _2300_;
  logic [31:0] _2301_;
  logic [31:0] _2302_;
  logic [15:0] _2303_;
  logic [31:0] _2304_;
  logic _2305_;
  logic [31:0] _2306_;
  logic [31:0] _2307_;
  logic [1:0] _2308_;
  logic [31:0] _2309_;
  logic _2310_;
  logic _2311_;
  logic _2312_;
  logic _2313_;
  logic [31:0] _2314_;
  logic _2315_;
  logic _2316_;
  logic _2317_;
  logic _2318_;
  logic _2319_;
  logic _2320_;
  logic _2321_;
  logic _2322_;
  logic _2323_;
  logic [31:0] _2324_;
  logic [31:0] _2325_;
  logic [31:0] _2326_;
  logic _2327_;
  logic [31:0] _2328_;
  logic [31:0] _2329_;
  logic [31:0] _2330_;
  logic [31:0] _2331_;
  logic [31:0] _2332_;
  logic [31:0] _2333_;
  logic [31:0] _2334_;
  logic [31:0] _2335_;
  logic _2336_;
  logic _2337_;
  logic _2338_;
  logic _2339_;
  logic _2340_;
  logic _2341_;
  logic _2342_;
  logic _2343_;
  logic _2344_;
  logic _2345_;
  logic _2346_;
  logic _2347_;
  logic _2348_;
  logic _2349_;
  logic _2350_;
  logic _2351_;
  logic _2352_;
  logic _2353_;
  logic _2354_;
  logic _2355_;
  logic _2356_;
  logic _2357_;
  logic _2358_;
  logic _2359_;
  logic _2360_;
  logic _2361_;
  logic _2362_;
  logic _2363_;
  logic _2364_;
  logic _2365_;
  logic _2366_;
  logic _2367_;
  logic _2368_;
  logic _2369_;
  logic _2370_;
  logic _2371_;
  logic _2372_;
  logic _2373_;
  logic _2374_;
  logic _2375_;
  logic _2376_;
  logic _2377_;
  logic _2378_;
  logic _2379_;
  logic _2380_;
  logic _2381_;
  logic _2382_;
  logic _2383_;
  logic _2384_;
  logic _2385_;
  logic _2386_;
  logic _2387_;
  logic _2388_;
  logic _2389_;
  logic _2390_;
  logic _2391_;
  logic _2392_;
  logic _2393_;
  logic _2394_;
  logic _2395_;
  logic _2396_;
  logic _2397_;
  logic _2398_;
  logic _2399_;
  logic _2400_;
  logic _2401_;
  logic _2402_;
  logic _2403_;
  logic _2404_;
  logic _2405_;
  logic _2406_;
  logic _2407_;
  logic _2408_;
  logic _2409_;
  logic _2410_;
  logic _2411_;
  logic _2412_;
  logic _2413_;
  logic _2414_;
  logic _2415_;
  logic _2416_;
  logic _2417_;
  logic _2418_;
  logic _2419_;
  logic _2420_;
  logic _2421_;
  logic _2422_;
  logic _2423_;
  logic _2424_;
  logic _2425_;
  logic _2426_;
  logic _2427_;
  logic _2428_;
  logic _2429_;
  logic _2430_;
  logic _2431_;
  logic _2432_;
  logic _2433_;
  logic _2434_;
  logic _2435_;
  logic _2436_;
  logic _2437_;
  logic _2438_;
  logic _2439_;
  logic _2440_;
  logic _2441_;
  logic _2442_;
  logic _2443_;
  logic _2444_;
  logic _2445_;
  logic _2446_;
  logic _2447_;
  logic _2448_;
  logic _2449_;
  logic _2450_;
  logic _2451_;
  logic _2452_;
  logic _2453_;
  logic _2454_;
  logic _2455_;
  logic _2456_;
  logic _2457_;
  logic _2458_;
  logic _2459_;
  logic _2460_;
  logic _2461_;
  logic _2462_;
  logic _2463_;
  logic _2464_;
  logic _2465_;
  logic _2466_;
  logic _2467_;
  logic _2468_;
  logic _2469_;
  logic _2470_;
  logic _2471_;
  logic _2472_;
  logic _2473_;
  logic _2474_;
  logic _2475_;
  logic _2476_;
  logic _2477_;
  logic _2478_;
  logic _2479_;
  logic _2480_;
  logic _2481_;
  logic _2482_;
  logic _2483_;
  logic _2484_;
  logic _2485_;
  logic _2486_;
  logic _2487_;
  logic _2488_;
  logic _2489_;
  logic _2490_;
  logic _2491_;
  logic _2492_;
  logic _2493_;
  logic _2494_;
  logic _2495_;
  logic _2496_;
  logic _2497_;
  logic _2498_;
  logic _2499_;
  logic _2500_;
  logic _2501_;
  logic _2502_;
  logic _2503_;
  logic _2504_;
  logic _2505_;
  logic _2506_;
  logic _2507_;
  logic _2508_;
  logic _2509_;
  logic _2510_;
  logic _2511_;
  logic _2512_;
  logic _2513_;
  logic _2514_;
  logic _2515_;
  logic _2516_;
  logic _2517_;
  logic _2518_;
  logic _2519_;
  logic _2520_;
  logic _2521_;
  logic _2522_;
  logic _2523_;
  logic _2524_;
  logic _2525_;
  logic _2526_;
  logic _2527_;
  logic _2528_;
  logic _2529_;
  logic _2530_;
  logic _2531_;
  logic _2532_;
  logic [31:0] _2533_;
  logic [31:0] _2534_;
  logic [31:0] _2535_;
  logic [31:0] _2536_;
  logic [31:0] _2537_;
  logic [31:0] _2538_;
  logic [31:0] _2539_;
  logic [31:0] _2540_;
  logic _2541_;
  logic _2542_;
  logic _2543_;
  logic _2544_;
  logic _2545_;
  logic _2546_;
  logic _2547_;
  logic _2548_;
  logic _2549_;
  logic _2550_;
  logic _2551_;
  logic _2552_;
  logic _2553_;
  logic _2554_;
  logic _2555_;
  logic _2556_;
  logic _2557_;
  logic _2558_;
  logic _2559_;
  logic _2560_;
  logic _2561_;
  logic _2562_;
  logic _2563_;
  logic _2564_;
  logic _2565_;
  logic _2566_;
  logic _2567_;
  logic _2568_;
  logic _2569_;
  logic _2570_;
  logic _2571_;
  logic _2572_;
  logic _2573_;
  logic _2574_;
  logic _2575_;
  logic _2576_;
  logic _2577_;
  logic _2578_;
  logic _2579_;
  logic _2580_;
  logic _2581_;
  logic _2582_;
  logic _2583_;
  logic _2584_;
  logic _2585_;
  logic _2586_;
  logic _2587_;
  logic _2588_;
  logic _2589_;
  logic _2590_;
  logic _2591_;
  logic _2592_;
  logic _2593_;
  logic _2594_;
  logic _2595_;
  logic _2596_;
  logic _2597_;
  logic _2598_;
  logic _2599_;
  logic _2600_;
  logic _2601_;
  logic _2602_;
  logic _2603_;
  logic _2604_;
  logic _2605_;
  logic _2606_;
  logic _2607_;
  logic _2608_;
  logic _2609_;
  logic _2610_;
  logic _2611_;
  logic _2612_;
  logic _2613_;
  logic _2614_;
  logic _2615_;
  logic _2616_;
  logic _2617_;
  logic _2618_;
  logic _2619_;
  logic _2620_;
  logic _2621_;
  logic _2622_;
  logic _2623_;
  logic _2624_;
  logic _2625_;
  logic _2626_;
  logic _2627_;
  logic _2628_;
  logic _2629_;
  logic _2630_;
  logic _2631_;
  logic _2632_;
  logic _2633_;
  logic _2634_;
  logic _2635_;
  logic _2636_;
  logic _2637_;
  logic _2638_;
  logic _2639_;
  logic _2640_;
  logic _2641_;
  logic _2642_;
  logic _2643_;
  logic _2644_;
  logic _2645_;
  logic _2646_;
  logic _2647_;
  logic _2648_;
  logic _2649_;
  logic _2650_;
  logic _2651_;
  logic _2652_;
  logic _2653_;
  logic _2654_;
  logic _2655_;
  logic _2656_;
  logic _2657_;
  logic _2658_;
  logic _2659_;
  logic _2660_;
  logic _2661_;
  logic _2662_;
  logic _2663_;
  logic _2664_;
  logic _2665_;
  logic _2666_;
  logic _2667_;
  logic _2668_;
  logic _2669_;
  logic _2670_;
  logic _2671_;
  logic _2672_;
  logic _2673_;
  logic _2674_;
  logic _2675_;
  logic _2676_;
  logic _2677_;
  logic _2678_;
  logic _2679_;
  logic _2680_;
  logic _2681_;
  logic _2682_;
  logic _2683_;
  logic _2684_;
  logic _2685_;
  logic _2686_;
  logic _2687_;
  logic _2688_;
  logic _2689_;
  logic _2690_;
  logic _2691_;
  logic _2692_;
  logic _2693_;
  logic _2694_;
  logic _2695_;
  logic _2696_;
  logic _2697_;
  logic _2698_;
  logic _2699_;
  logic _2700_;
  logic _2701_;
  logic _2702_;
  logic _2703_;
  logic _2704_;
  logic _2705_;
  logic _2706_;
  logic _2707_;
  logic _2708_;
  logic _2709_;
  logic _2710_;
  logic _2711_;
  logic _2712_;
  logic _2713_;
  logic _2714_;
  logic _2715_;
  logic _2716_;
  logic _2717_;
  logic _2718_;
  logic _2719_;
  logic _2720_;
  logic _2721_;
  logic _2722_;
  logic _2723_;
  logic _2724_;
  logic _2725_;
  logic _2726_;
  logic _2727_;
  logic _2728_;
  logic _2729_;
  logic _2730_;
  logic _2731_;
  logic _2732_;
  logic _2733_;
  logic _2734_;
  logic _2735_;
  logic _2736_;
  logic _2737_;
  logic [2:0] _2738_;
  logic [1:0] _2739_;
  logic [1:0] _2740_;
  logic [1:0] _2741_;
  logic _2742_;
  logic _2743_;
  logic _2744_;
  logic [1:0] _2745_;
  logic _2746_;
  logic _2747_;
  logic _2748_;
  logic [31:0] _2749_;
  logic [31:0] _2750_;
  logic _2751_;
  logic _2752_;
  logic _2753_;
  logic _2754_;
  logic _2755_;
  logic _2756_;
  logic _2757_;
  logic _2758_;
  logic _2759_;
  logic _2760_;
  logic _2761_;
  logic _2762_;
  logic _2763_;
  logic [1:0] _2764_;
  logic [63:0] _2765_;
  logic [63:0] _2766_;
  logic _2767_;
  logic _2768_;
  logic _2769_;
  logic _2770_;
  logic [1:0] _2771_;
  logic [1:0] _2772_;
  logic [1:0] _2773_;
  logic _2774_;
  logic _2775_;
  logic _2776_;
  logic _2777_;
  logic [31:0] _2778_;
  logic _2779_;
  logic [31:0] _2780_;
  logic _2781_;
  logic _2782_;
  logic [31:0] _2783_;
  logic [31:0] _2784_;
  logic [1:0] _2785_;
  logic [99:0] _2786_;
  logic _2787_;
  logic _2788_;
  logic _2789_;
  logic _2790_;
  logic _2791_;
  logic _2792_;
  logic _2793_;
  logic _2794_;
  logic _2795_;
  logic _2796_;
  logic _2797_;
  logic _2798_;
  logic _2799_;
  logic _2800_;
  logic _2801_;
  logic _2802_;
  logic _2803_;
  logic _2804_;
  logic _2805_;
  logic _2806_;
  logic _2807_;
  logic _2808_;
  logic _2809_;
  logic _2810_;
  logic [31:0] _2811_;
  logic [31:0] _2812_;
  logic _2813_;
  logic _2814_;
  logic _2815_;
  logic [99:0] _2816_;
  logic [1:0] _2817_;
  logic [1:0] _2818_;
  logic [31:0] _2819_;
  logic [31:0] _2820_;
  logic [31:0] _2821_;
  logic [31:0] _2822_;
  logic _2823_;
  logic _2824_;
  logic _2825_;
  logic _2826_;
  logic [1:0] _2827_;
  logic [1:0] _2828_;
  logic [1:0] _2829_;
  logic [1:0] _2830_;
  logic [1:0] _2831_;
  logic _2832_;
  logic _2833_;
  logic [31:0] _2834_;
  logic [31:0] _2835_;
  logic [31:0] _2836_;
  logic [31:0] _2837_;
  logic [31:0] _2838_;
  logic [2:0] _2839_;
  logic [2:0] _2840_;
  logic _2841_;
  logic _2842_;
  logic _2843_;
  logic [31:0] _2844_;
  logic _2845_;
  logic _2846_;
  logic _2847_;
  logic _2848_;
  logic _2849_;
  logic [31:0] _2850_;
  logic _2851_;
  logic _2852_;
  logic _2853_;
  logic _2854_;
  logic _2855_;
  logic [31:0] _2856_;
  logic _2857_;
  logic _2858_;
  logic _2859_;
  logic _2860_;
  logic _2861_;
  logic [31:0] _2862_;
  logic _2863_;
  logic _2864_;
  logic _2865_;
  logic _2866_;
  logic _2867_;
  logic [31:0] _2868_;
  logic _2869_;
  logic _2870_;
  logic _2871_;
  logic _2872_;
  logic _2873_;
  logic [31:0] _2874_;
  logic _2875_;
  logic _2876_;
  logic _2877_;
  logic _2878_;
  logic _2879_;
  logic [31:0] _2880_;
  logic _2881_;
  logic _2882_;
  logic _2883_;
  logic _2884_;
  logic _2885_;
  logic [31:0] _2886_;
  logic _2887_;
  logic _2888_;
  logic _2889_;
  logic _2890_;
  logic _2891_;
  logic [31:0] _2892_;
  logic _2893_;
  logic _2894_;
  logic _2895_;
  logic _2896_;
  logic _2897_;
  logic _2898_;
  logic [31:0] _2899_;
  logic _2900_;
  logic _2901_;
  logic [2:0] _2902_;
  logic [2:0] _2903_;
  logic _2904_;
  logic _2905_;
  logic _2906_;
  logic _2907_;
  logic [31:0] _2908_;
  logic _2909_;
  logic _2910_;
  logic _2911_;
  logic [2:0] _2912_;
  logic _2913_;
  logic _2914_;
  logic _2915_;
  logic _2916_;
  logic [31:0] _2917_;
  logic _2918_;
  logic _2919_;
  logic [1:0] _2920_;
  logic [2:0] _2921_;
  logic _2922_;
  logic _2923_;
  logic _2924_;
  logic _2925_;
  logic [31:0] _2926_;
  logic _2927_;
  logic _2928_;
  logic [1:0] _2929_;
  logic _2930_;
  logic _2931_;
  logic _2932_;
  logic _2933_;
  logic [31:0] _2934_;
  logic _2935_;
  logic _2936_;
  logic [2:0] _2937_;
  logic _2938_;
  logic _2939_;
  logic _2940_;
  logic _2941_;
  logic [31:0] _2942_;
  logic _2943_;
  logic _2944_;
  logic [2:0] _2945_;
  logic _2946_;
  logic _2947_;
  logic _2948_;
  logic _2949_;
  logic [31:0] _2950_;
  logic _2951_;
  logic _2952_;
  logic [2:0] _2953_;
  logic _2954_;
  logic [2:0] _2955_;
  logic [2:0] _2956_;
  logic [31:0] _2957_;
  logic [31:0] _2958_;
  logic _2959_;
  logic _2960_;
  logic _2961_;
  logic _2962_;
  logic _2963_;
  logic _2964_;
  logic _2965_;
  logic [31:0] _2966_;
  logic [31:0] _2967_;
  logic _2968_;
  logic _2969_;
  logic _2970_;
  logic _2971_;
  logic _2972_;
  logic _2973_;
  logic _2974_;
  logic _2975_;
  logic _2976_;
  logic _2977_;
  logic _2978_;
  logic _2979_;
  logic _2980_;
  logic _2981_;
  logic _2982_;
  logic _2983_;
  logic _2984_;
  logic _2985_;
  logic _2986_;
  logic _2987_;
  logic _2988_;
  logic _2989_;
  logic _2990_;
  logic _2991_;
  logic _2992_;
  logic _2993_;
  logic _2994_;
  logic _2995_;
  logic _2996_;
  logic _2997_;
  logic _2998_;
  logic [1:0] _2999_;
  logic [1:0] _3000_;
  logic _3001_;
  logic _3002_;
  logic _3003_;
  logic _3004_;
  logic _3005_;
  logic _3006_;
  logic _3007_;
  logic _3008_;
  logic _3009_;
  logic _3010_;
  logic _3011_;
  logic _3012_;
  logic _3013_;
  logic _3014_;
  logic _3015_;
  logic _3016_;
  logic _3017_;
  logic _3018_;
  logic _3019_;
  logic _3020_;
  logic _3021_;
  logic _3022_;
  logic _3023_;
  logic _3024_;
  logic [31:0] _3025_;
  logic [31:0] _3026_;
  logic [31:0] _3027_;
  logic [31:0] _3028_;
  logic [31:0] _3029_;
  logic [31:0] _3030_;
  logic [31:0] _3031_;
  logic [31:0] _3032_;
  logic [31:0] _3033_;
  logic [31:0] _3034_;
  logic [31:0] _3035_;
  logic [31:0] _3036_;
  logic [31:0] _3037_;
  logic [31:0] _3038_;
  logic [31:0] _3039_;
  logic [31:0] _3040_;
  logic _3041_;
  logic _3042_;
  logic _3043_;
  logic _3044_;
  logic [31:0] _3045_;
  logic _3046_;
  logic _3047_;
  logic _3048_;
  logic [31:0] _3049_;
  logic [31:0] _3050_;
  logic [31:0] _3051_;
  logic [31:0] _3052_;
  logic [31:0] _3053_;
  logic [1:0] _3054_;
  logic [1:0] _3055_;
  logic [1:0] _3056_;
  logic [31:0] _3057_;
  logic [31:0] _3058_;
  logic [31:0] _3059_;
  logic [2:0] _3060_;
  logic [2:0] _3061_;
  logic [2:0] _3062_;
  logic [31:0] _3063_;
  logic [31:0] _3064_;
  logic [31:0] _3065_;
  logic [1:0] _3066_;
  logic [15:0] _3067_;
  logic [15:0] _3068_;
  logic [15:0] _3069_;
  logic [15:0] _3070_;
  logic _3071_;
  logic _3072_;
  logic [31:0] _3073_;
  logic [31:0] _3074_;
  logic [31:0] _3075_;
  logic [31:0] _3076_;
  logic [31:0] _3077_;
  logic [31:0] _3078_;
  logic [31:0] _3079_;
  logic [31:0] _3080_;
  logic [31:0] _3081_;
  logic [31:0] _3082_;
  logic _3083_;
  logic _3084_;
  logic [1:0] _3085_;
  logic [31:0] _3086_;
  logic [31:0] _3087_;
  logic _3088_;
  logic _3089_;
  logic _3090_;
  logic _3091_;
  logic [31:0] _3092_;
  logic _3093_;
  logic _3094_;
  logic [31:0] _3095_;
  logic [31:0] _3096_;
  logic [31:0] _3097_;
  logic [31:0] _3098_;
  logic _3099_;
  logic [31:0] _3100_;
  logic _3101_;
  logic [31:0] _3102_;
  logic [31:0] _3103_;
  logic [31:0] _3104_;
  logic [31:0] _3105_;
  logic _3106_;
  logic [31:0] _3107_;
  logic [31:0] _3108_;
  logic [31:0] _3109_;
  logic [31:0] _3110_;
  logic [31:0] _3111_;
  logic [31:0] _3112_;
  logic [31:0] _3113_;
  logic [31:0] _3114_;
  logic [31:0] _3115_;
  logic [31:0] _3116_;
  logic [31:0] _3117_;
  logic [31:0] _3118_;
  logic [31:0] _3119_;
  logic [31:0] _3120_;
  logic [31:0] _3121_;
  logic [31:0] _3122_;
  logic _3123_;
  logic _3124_;
  logic _3125_;
  logic _3126_;
  logic _3127_;
  logic _3128_;
  logic _3129_;
  logic _3130_;
  logic _3131_;
  logic _3132_;
  logic _3133_;
  logic _3134_;
  logic _3135_;
  logic _3136_;
  logic _3137_;
  logic _3138_;
  logic _3139_;
  logic _3140_;
  logic _3141_;
  logic _3142_;
  logic _3143_;
  logic _3144_;
  logic _3145_;
  logic _3146_;
  logic _3147_;
  logic _3148_;
  logic _3149_;
  logic _3150_;
  logic _3151_;
  logic _3152_;
  logic _3153_;
  logic _3154_;
  logic _3155_;
  logic _3156_;
  logic _3157_;
  logic _3158_;
  logic _3159_;
  logic _3160_;
  logic _3161_;
  logic _3162_;
  logic _3163_;
  logic _3164_;
  logic _3165_;
  logic _3166_;
  logic _3167_;
  logic _3168_;
  logic _3169_;
  logic _3170_;
  logic _3171_;
  logic _3172_;
  logic _3173_;
  logic _3174_;
  logic _3175_;
  logic _3176_;
  logic _3177_;
  logic _3178_;
  logic _3179_;
  logic _3180_;
  logic _3181_;
  logic _3182_;
  logic _3183_;
  logic _3184_;
  logic _3185_;
  logic _3186_;
  logic _3187_;
  logic _3188_;
  logic _3189_;
  logic _3190_;
  logic _3191_;
  logic _3192_;
  logic _3193_;
  logic _3194_;
  logic _3195_;
  logic _3196_;
  logic _3197_;
  logic _3198_;
  logic _3199_;
  logic _3200_;
  logic _3201_;
  logic _3202_;
  logic _3203_;
  logic _3204_;
  logic _3205_;
  logic _3206_;
  logic _3207_;
  logic _3208_;
  logic _3209_;
  logic _3210_;
  logic _3211_;
  logic _3212_;
  logic _3213_;
  logic _3214_;
  logic _3215_;
  logic _3216_;
  logic _3217_;
  logic _3218_;
  logic _3219_;
  logic _3220_;
  logic _3221_;
  logic _3222_;
  logic _3223_;
  logic _3224_;
  logic _3225_;
  logic _3226_;
  logic _3227_;
  logic _3228_;
  logic _3229_;
  logic _3230_;
  logic _3231_;
  logic _3232_;
  logic [5:0] _3233_;
  logic [5:0] _3234_;
  logic _3235_;
  logic _3236_;
  logic _3237_;
  logic _3238_;
  logic _3239_;
  logic _3240_;
  logic _3241_;
  logic _3242_;
  logic _3243_;
  logic _3244_;
  logic _3245_;
  logic _3246_;
  logic _3247_;
  logic _3248_;
  logic _3249_;
  logic _3250_;
  logic _3251_;
  logic _3252_;
  logic _3253_;
  logic _3254_;
  logic _3255_;
  logic _3256_;
  logic _3257_;
  logic _3258_;
  logic _3259_;
  logic _3260_;
  logic _3261_;
  logic _3262_;
  logic _3263_;
  logic _3264_;
  logic _3265_;
  logic _3266_;
  logic _3267_;
  logic _3268_;
  logic _3269_;
  logic _3270_;
  logic _3271_;
  logic _3272_;
  logic _3273_;
  logic _3274_;
  logic _3275_;
  logic _3276_;
  logic _3277_;
  logic _3278_;
  logic _3279_;
  logic _3280_;
  logic _3281_;
  logic _3282_;
  logic _3283_;
  logic _3284_;
  logic _3285_;
  logic _3286_;
  logic _3287_;
  logic _3288_;
  logic _3289_;
  logic _3290_;
  logic _3291_;
  logic _3292_;
  logic _3293_;
  logic _3294_;
  logic _3295_;
  logic _3296_;
  logic _3297_;
  logic _3298_;
  logic _3299_;
  logic _3300_;
  logic _3301_;
  logic _3302_;
  logic _3303_;
  logic _3304_;
  logic _3305_;
  logic _3306_;
  logic _3307_;
  logic _3308_;
  logic _3309_;
  logic _3310_;
  logic _3311_;
  logic _3312_;
  logic _3313_;
  logic _3314_;
  logic _3315_;
  logic _3316_;
  logic _3317_;
  logic _3318_;
  logic _3319_;
  logic _3320_;
  logic _3321_;
  logic _3322_;
  logic _3323_;
  logic _3324_;
  logic _3325_;
  logic _3326_;
  logic _3327_;
  logic _3328_;
  logic _3329_;
  logic _3330_;
  logic _3331_;
  logic _3332_;
  logic _3333_;
  logic _3334_;
  logic _3335_;
  logic _3336_;
  logic _3337_;
  logic _3338_;
  logic _3339_;
  logic _3340_;
  logic _3341_;
  logic _3342_;
  logic _3343_;
  logic _3344_;
  logic _3345_;
  logic _3346_;
  logic _3347_;
  logic _3348_;
  logic _3349_;
  logic _3350_;
  logic _3351_;
  logic _3352_;
  logic _3353_;
  logic _3354_;
  logic _3355_;
  logic _3356_;
  logic _3357_;
  logic _3358_;
  logic _3359_;
  logic _3360_;
  logic _3361_;
  logic _3362_;
  logic _3363_;
  logic _3364_;
  logic _3365_;
  logic _3366_;
  logic _3367_;
  logic _3368_;
  logic _3369_;
  logic _3370_;
  logic _3371_;
  logic _3372_;
  logic _3373_;
  logic _3374_;
  logic _3375_;
  logic _3376_;
  logic _3377_;
  logic _3378_;
  logic _3379_;
  logic _3380_;
  logic _3381_;
  logic _3382_;
  logic _3383_;
  logic _3384_;
  logic _3385_;
  logic _3386_;
  logic _3387_;
  logic _3388_;
  logic _3389_;
  logic _3390_;
  logic _3391_;
  logic _3392_;
  logic _3393_;
  logic _3394_;
  logic _3395_;
  logic _3396_;
  logic _3397_;
  logic _3398_;
  logic _3399_;
  logic _3400_;
  logic _3401_;
  logic _3402_;
  logic _3403_;
  logic _3404_;
  logic _3405_;
  logic _3406_;
  logic _3407_;
  logic _3408_;
  logic _3409_;
  logic _3410_;
  logic _3411_;
  logic [31:0] _3412_;
  logic [31:0] _3413_;
  logic [31:0] _3414_;
  logic [31:0] _3415_;
  logic [31:0] _3416_;
  logic _3417_;
  logic _3418_;
  logic _3419_;
  logic _3420_;
  logic _3421_;
  logic _3422_;
  logic _3423_;
  logic _3424_;
  logic _3425_;
  logic [31:0] _3426_;
  logic [31:0] _3427_;
  logic _3428_;
  logic _3429_;
  logic [9:0] _3430_;
  logic [9:0] _3431_;
  logic [9:0] _3432_;
  logic [5:0] _3433_;
  logic [5:0] _3434_;
  logic [5:0] _3435_;
  logic [31:0] _3436_;
  logic [31:0] _3437_;
  logic [31:0] _3438_;
  logic [31:0] _3439_;
  logic [31:0] _3440_;
  logic [31:0] _3441_;
  logic [31:0] _3442_;
  logic [31:0] _3443_;
  logic _3444_;
  logic _3445_;
  logic _3446_;
  logic _3447_;
  logic [31:0] _3448_;
  logic _3449_;
  logic _3450_;
  logic _3451_;
  logic _3452_;
  logic _3453_;
  logic _3454_;
  logic _3455_;
  logic _3456_;
  logic _3457_;
  logic _3458_;
  logic [9:0] _3459_;
  logic [5:0] _3460_;
  logic _3461_;
  logic _3462_;
  logic _3463_;
  logic _3464_;
  logic _3465_;
  logic _3466_;
  logic _3467_;
  logic _3468_;
  logic _3469_;
  logic _3470_;
  logic _3471_;
  logic _3472_;
  logic _3473_;
  logic _3474_;
  logic _3475_;
  logic _3476_;
  logic _3477_;
  logic _3478_;
  logic _3479_;
  logic _3480_;
  logic _3481_;
  logic _3482_;
  logic _3483_;
  logic _3484_;
  logic _3485_;
  logic _3486_;
  logic _3487_;
  logic _3488_;
  logic _3489_;
  logic [5:0] _3490_;
  logic [5:0] _3491_;
  logic [31:0] _3492_;
  logic [31:0] _3493_;
  logic [31:0] _3494_;
  logic [31:0] _3495_;
  logic [31:0] _3496_;
  logic [31:0] _3497_;
  logic [31:0] _3498_;
  logic [31:0] _3499_;
  logic [31:0] _3500_;
  logic [31:0] _3501_;
  logic _3502_;
  logic _3503_;
  logic [9:0] _3504_;
  logic [9:0] _3505_;
  logic [9:0] _3506_;
  logic _3507_;
  logic [5:0] _3508_;
  logic _3509_;
  logic _3510_;
  logic _3511_;
  logic _3512_;
  logic [5:0] _3513_;
  logic _3514_;
  logic [5:0] _3515_;
  logic [5:0] _3516_;
  logic [5:0] _3517_;
  logic [31:0] _3518_;
  logic [31:0] _3519_;
  logic [31:0] _3520_;
  logic [31:0] _3521_;
  logic [31:0] _3522_;
  logic [31:0] _3523_;
  logic _3524_;
  logic _3525_;
  logic [9:0] _3526_;
  logic [9:0] _3527_;
  logic _3528_;
  logic _3529_;
  logic _3530_;
  logic _3531_;
  logic [31:0] _3532_;
  logic [31:0] _3533_;
  logic [31:0] _3534_;
  logic [31:0] _3535_;
  logic _3536_;
  logic _3537_;
  logic _3538_;
  logic _3539_;
  logic _3540_;
  logic _3541_;
  logic _3542_;
  logic _3543_;
  logic _3544_;
  logic _3545_;
  logic _3546_;
  logic _3547_;
  logic _3548_;
  logic _3549_;
  logic _3550_;
  logic _3551_;
  logic _3552_;
  logic _3553_;
  logic _3554_;
  logic _3555_;
  logic [31:0] _3556_;
  logic [31:0] _3557_;
  logic [31:0] _3558_;
  logic [31:0] _3559_;
  logic _3560_;
  logic [5:0] _3561_;
  logic [5:0] _3562_;
  logic _3563_;
  logic [5:0] _3564_;
  logic [9:0] _3565_;
  logic [9:0] _3566_;
  logic [9:0] _3567_;
  logic [5:0] _3568_;
  logic [5:0] _3569_;
  logic [5:0] _3570_;
  logic [31:0] _3571_;
  logic [31:0] _3572_;
  logic [31:0] _3573_;
  logic [31:0] _3574_;
  logic [31:0] _3575_;
  logic [31:0] _3576_;
  logic [31:0] _3577_;
  logic [31:0] _3578_;
  logic _3579_;
  logic _3580_;
  logic _3581_;
  logic _3582_;
  logic [31:0] _3583_;
  logic _3584_;
  logic _3585_;
  logic _3586_;
  logic _3587_;
  logic _3588_;
  logic _3589_;
  logic _3590_;
  logic _3591_;
  logic _3592_;
  logic _3593_;
  logic [9:0] _3594_;
  logic [5:0] _3595_;
  logic _3596_;
  logic _3597_;
  logic _3598_;
  logic _3599_;
  logic _3600_;
  logic _3601_;
  logic _3602_;
  logic _3603_;
  logic _3604_;
  logic _3605_;
  logic _3606_;
  logic _3607_;
  logic _3608_;
  logic _3609_;
  logic _3610_;
  logic _3611_;
  logic _3612_;
  logic _3613_;
  logic _3614_;
  logic _3615_;
  logic _3616_;
  logic _3617_;
  logic _3618_;
  logic _3619_;
  logic _3620_;
  logic _3621_;
  logic _3622_;
  logic _3623_;
  logic _3624_;
  logic [5:0] _3625_;
  logic [5:0] _3626_;
  logic [31:0] _3627_;
  logic [31:0] _3628_;
  logic [31:0] _3629_;
  logic [31:0] _3630_;
  logic [31:0] _3631_;
  logic [31:0] _3632_;
  logic [31:0] _3633_;
  logic [31:0] _3634_;
  logic [9:0] _3635_;
  logic [9:0] _3636_;
  logic [9:0] _3637_;
  logic _3638_;
  logic [5:0] _3639_;
  logic _3640_;
  logic _3641_;
  logic _3642_;
  logic _3643_;
  logic [5:0] _3644_;
  logic _3645_;
  logic [5:0] _3646_;
  logic [5:0] _3647_;
  logic [5:0] _3648_;
  logic [31:0] _3649_;
  logic [31:0] _3650_;
  logic [31:0] _3651_;
  logic [31:0] _3652_;
  logic [9:0] _3653_;
  logic [9:0] _3654_;
  logic _3655_;
  logic _3656_;
  logic _3657_;
  logic _3658_;
  logic [31:0] _3659_;
  logic [31:0] _3660_;
  logic [31:0] _3661_;
  logic [31:0] _3662_;
  logic _3663_;
  logic _3664_;
  logic _3665_;
  logic _3666_;
  logic _3667_;
  logic _3668_;
  logic _3669_;
  logic _3670_;
  logic _3671_;
  logic _3672_;
  logic _3673_;
  logic _3674_;
  logic _3675_;
  logic _3676_;
  logic _3677_;
  logic _3678_;
  logic _3679_;
  logic _3680_;
  logic _3681_;
  logic _3682_;
  logic [31:0] _3683_;
  logic [31:0] _3684_;
  logic [31:0] _3685_;
  logic [31:0] _3686_;
  logic _3687_;
  logic [5:0] _3688_;
  logic [5:0] _3689_;
  logic _3690_;
  logic [5:0] _3691_;
  logic [31:0] _3692_;
  logic [31:0] _3693_;
  logic [31:0] _3694_;
  logic [31:0] _3695_;
  logic [31:0] _3696_;
  logic [31:0] _3697_;
  logic [31:0] _3698_;
  logic [31:0] _3699_;
  logic [31:0] _3700_;
  logic [31:0] _3701_;
  logic [31:0] _3702_;
  logic [31:0] _3703_;
  logic [31:0] _3704_;
  logic [31:0] _3705_;
  logic [31:0] _3706_;
  logic [31:0] _3707_;
  logic [31:0] _3708_;
  logic [31:0] _3709_;
  logic [31:0] _3710_;
  logic [31:0] _3711_;
  logic [31:0] _3712_;
  logic [31:0] _3713_;
  logic [31:0] _3714_;
  logic [31:0] _3715_;
  logic [31:0] _3716_;
  logic [31:0] _3717_;
  logic [31:0] _3718_;
  logic [31:0] _3719_;
  logic [31:0] _3720_;
  logic [31:0] _3721_;
  logic [31:0] _3722_;
  logic _3723_;
  logic _3724_;
  logic _3725_;
  logic _3726_;
  logic _3727_;
  logic _3728_;
  logic _3729_;
  logic _3730_;
  logic _3731_;
  logic _3732_;
  logic _3733_;
  logic _3734_;
  logic _3735_;
  logic _3736_;
  logic _3737_;
  logic _3738_;
  logic _3739_;
  logic _3740_;
  logic _3741_;
  logic _3742_;
  logic _3743_;
  logic _3744_;
  logic _3745_;
  logic _3746_;
  logic _3747_;
  logic _3748_;
  logic _3749_;
  logic _3750_;
  logic _3751_;
  logic _3752_;
  logic _3753_;
  logic _3754_;
  logic _3755_;
  logic _3756_;
  logic _3757_;
  logic _3758_;
  logic _3759_;
  logic _3760_;
  logic _3761_;
  logic _3762_;
  logic _3763_;
  logic _3764_;
  logic _3765_;
  logic _3766_;
  logic _3767_;
  logic _3768_;
  logic _3769_;
  logic _3770_;
  logic _3771_;
  logic _3772_;
  logic _3773_;
  logic _3774_;
  logic _3775_;
  logic _3776_;
  logic _3777_;
  logic _3778_;
  logic _3779_;
  logic _3780_;
  logic _3781_;
  logic _3782_;
  logic _3783_;
  logic _3784_;
  logic _3785_;
  logic _3786_;
  logic _3787_;
  logic _3788_;
  logic _3789_;
  logic _3790_;
  logic _3791_;
  logic _3792_;
  logic _3793_;
  logic _3794_;
  logic _3795_;
  logic _3796_;
  logic _3797_;
  logic _3798_;
  logic _3799_;
  logic _3800_;
  logic _3801_;
  logic _3802_;
  logic _3803_;
  logic _3804_;
  logic _3805_;
  logic _3806_;
  logic _3807_;
  logic _3808_;
  logic _3809_;
  logic _3810_;
  logic _3811_;
  logic _3812_;
  logic _3813_;
  logic _3814_;
  logic _3815_;
  logic _3816_;
  logic _3817_;
  logic _3818_;
  logic _3819_;
  logic _3820_;
  logic _3821_;
  logic _3822_;
  logic _3823_;
  logic _3824_;
  logic _3825_;
  logic _3826_;
  logic _3827_;
  logic _3828_;
  logic _3829_;
  logic _3830_;
  logic _3831_;
  logic _3832_;
  logic _3833_;
  logic _3834_;
  logic _3835_;
  logic _3836_;
  logic _3837_;
  logic _3838_;
  logic _3839_;
  logic _3840_;
  logic _3841_;
  logic _3842_;
  logic _3843_;
  logic _3844_;
  logic _3845_;
  logic _3846_;
  logic _3847_;
  logic _3848_;
  logic _3849_;
  logic _3850_;
  logic _3851_;
  logic _3852_;
  logic _3853_;
  logic _3854_;
  logic _3855_;
  logic _3856_;
  logic _3857_;
  logic _3858_;
  logic _3859_;
  logic _3860_;
  logic _3861_;
  logic _3862_;
  logic _3863_;
  logic _3864_;
  logic _3865_;
  logic _3866_;
  logic _3867_;
  logic _3868_;
  logic _3869_;
  logic _3870_;
  logic _3871_;
  logic _3872_;
  logic _3873_;
  logic _3874_;
  logic _3875_;
  logic _3876_;
  logic _3877_;
  logic _3878_;
  logic _3879_;
  logic _3880_;
  logic _3881_;
  logic _3882_;
  logic _3883_;
  logic _3884_;
  logic _3885_;
  logic _3886_;
  logic _3887_;
  logic _3888_;
  logic _3889_;
  logic _3890_;
  logic _3891_;
  logic _3892_;
  logic _3893_;
  logic _3894_;
  logic _3895_;
  logic _3896_;
  logic _3897_;
  logic _3898_;
  logic _3899_;
  logic _3900_;
  logic _3901_;
  logic _3902_;
  logic _3903_;
  logic _3904_;
  logic _3905_;
  logic _3906_;
  logic _3907_;
  logic _3908_;
  logic [31:0] _3909_;
  logic [31:0] _3910_;
  logic [31:0] _3911_;
  logic [31:0] _3912_;
  logic [31:0] _3913_;
  logic [31:0] _3914_;
  logic [31:0] _3915_;
  logic [31:0] _3916_;
  logic [31:0] _3917_;
  logic [31:0] _3918_;
  logic [31:0] _3919_;
  logic [31:0] _3920_;
  logic [31:0] _3921_;
  logic [31:0] _3922_;
  logic [31:0] _3923_;
  logic [31:0] _3924_;
  logic [31:0] _3925_;
  logic [31:0] _3926_;
  logic [31:0] _3927_;
  logic [31:0] _3928_;
  logic [31:0] _3929_;
  logic [31:0] _3930_;
  logic [31:0] _3931_;
  logic [31:0] _3932_;
  logic [31:0] _3933_;
  logic [31:0] _3934_;
  logic [31:0] _3935_;
  logic [31:0] _3936_;
  logic [31:0] _3937_;
  logic [31:0] _3938_;
  logic [31:0] _3939_;
  logic [31:0] _3940_;
  logic [31:0] _3941_;
  logic [31:0] _3942_;
  logic [31:0] _3943_;
  logic [31:0] _3944_;
  logic [31:0] _3945_;
  logic [31:0] _3946_;
  logic [31:0] _3947_;
  logic [31:0] _3948_;
  logic [31:0] _3949_;
  logic [31:0] _3950_;
  logic [31:0] _3951_;
  logic [31:0] _3952_;
  logic [31:0] _3953_;
  logic [31:0] _3954_;
  logic [31:0] _3955_;
  logic [31:0] _3956_;
  logic [31:0] _3957_;
  logic [31:0] _3958_;
  logic [31:0] _3959_;
  logic [31:0] _3960_;
  logic [31:0] _3961_;
  logic [31:0] _3962_;
  logic [31:0] _3963_;
  logic [31:0] _3964_;
  logic [31:0] _3965_;
  logic [31:0] _3966_;
  logic [31:0] _3967_;
  logic [31:0] _3968_;
  logic [31:0] _3969_;
  logic [31:0] _3970_;
  logic [31:0] _3971_;
  logic _3972_;
  logic [31:0] _3973_;
  logic _3974_;
  logic _3975_;
  logic _3976_;
  logic _3977_;
  logic _3978_;
  logic _3979_;
  logic _3980_;
  logic [3:0] _3981_;
  logic _3982_;
  logic _3983_;
  logic _3984_;
  logic _3985_;
  logic [31:0] _3986_;
  logic [31:0] _3987_;
  logic _3988_;
  logic [3:0] _3989_;
  logic [31:0] _3990_;
  logic [31:0] _3991_;
  logic [3:0] _3992_;
  logic [31:0] _3993_;
  logic [31:0] _3994_;
  logic [3:0] _3995_;
  logic [7:0] _3996_;
  logic [31:0] _3997_;
  logic [3:0] _3998_;
  logic [31:0] _3999_;
  logic [31:0] _4000_;
  logic [15:0] _4001_;
  logic [31:0] _4002_;
  logic [31:0] _4003_;
  logic [31:0] _4004_;
  logic _4005_;
  logic [31:0] _4006_;
  logic _4007_;
  logic _4008_;
  logic _4009_;
  logic [5:0] _4010_;
  logic [5:0] _4011_;
  logic [5:0] _4012_;
  logic _4013_;
  logic _4014_;
  logic _4015_;
  logic _4016_;
  logic _4017_;
  logic _4018_;
  logic _4019_;
  logic _4020_;
  logic _4021_;
  logic _4022_;
  logic _4023_;
  logic _4024_;
  logic _4025_;
  logic _4026_;
  logic _4027_;
  logic _4028_;
  logic _4029_;
  logic _4030_;
  logic _4031_;
  logic _4032_;
  logic _4033_;
  logic _4034_;
  logic _4035_;
  logic _4036_;
  logic _4037_;
  logic _4038_;
  logic _4039_;
  logic _4040_;
  logic _4041_;
  logic _4042_;
  logic _4043_;
  logic _4044_;
  logic _4045_;
  logic _4046_;
  logic _4047_;
  logic _4048_;
  logic _4049_;
  logic _4050_;
  logic _4051_;
  logic _4052_;
  logic _4053_;
  logic _4054_;
  logic _4055_;
  logic _4056_;
  logic _4057_;
  logic _4058_;
  logic _4059_;
  logic _4060_;
  logic _4061_;
  logic _4062_;
  logic _4063_;
  logic _4064_;
  logic _4065_;
  logic _4066_;
  logic _4067_;
  logic _4068_;
  logic _4069_;
  logic _4070_;
  logic _4071_;
  logic _4072_;
  logic [3:0] _4073_;
  logic _4074_;
  logic _4075_;
  logic _4076_;
  logic _4077_;
  logic _4078_;
  logic _4079_;
  logic _4080_;
  logic _4081_;
  logic _4082_;
  logic _4083_;
  logic _4084_;
  logic _4085_;
  logic _4086_;
  logic _4087_;
  logic _4088_;
  logic _4089_;
  logic _4090_;
  logic _4091_;
  logic _4092_;
  logic _4093_;
  logic _4094_;
  logic _4095_;
  logic _4096_;
  logic _4097_;
  logic _4098_;
  logic _4099_;
  logic _4100_;
  logic _4101_;
  logic _4102_;
  logic _4103_;
  logic _4104_;
  logic _4105_;
  logic _4106_;
  logic _4107_;
  logic [3:0] _4108_;
  logic [3:0] _4109_;
  logic [3:0] _4110_;
  logic _4111_;
  logic _4112_;
  logic _4113_;
  logic [31:0] _4114_;
  logic [31:0] _4115_;
  logic [31:0] _4116_;
  logic [31:0] _4117_;
  logic [31:0] _4118_;
  logic [31:0] _4119_;
  logic _4120_;
  logic _4121_;
  logic _4122_;
  logic _4123_;
  logic _4124_;
  logic _4125_;
  logic _4126_;
  logic _4127_;
  logic [5:0] _4128_;
  logic [5:0] _4129_;
  logic [35:0] _4130_;
  logic [35:0] _4131_;
  logic [1:0] _4132_;
  logic _4133_;
  logic _4134_;
  logic _4135_;
  logic [31:0] _4136_;
  logic [1:0] _4137_;
  logic _4138_;
  logic _4139_;
  logic _4140_;
  logic _4141_;
  logic _4142_;
  logic _4143_;
  logic [35:0] _4144_;
  logic [1:0] _4145_;
  logic [1:0] _4146_;
  logic _4147_;
  logic _4148_;
  logic [31:0] _4149_;
  logic _4150_;
  logic [32:0] _4151_;
  logic [32:0] _4152_;
  logic [31:0] _4153_;
  logic [32:0] _4154_;
  logic [32:0] _4155_;
  logic [31:0] _4156_;
  logic _4157_;
  logic _4158_;
  logic _4159_;
  logic _4160_;
  logic _4161_;
  logic _4162_;
  logic _4163_;
  logic _4164_;
  logic [31:0] _4165_;
  logic _4166_;
  logic _4167_;
  logic [32:0] _4168_;
  logic [32:0] _4169_;
  logic [32:0] _4170_;
  logic [32:0] _4171_;
  logic [31:0] branch_csr_pc_w;
  logic branch_csr_request_w;
  logic [31:0] branch_d_exec0_pc_w;
  logic branch_d_exec0_request_w;
  logic [31:0] branch_d_exec1_pc_w;
  logic branch_d_exec1_request_w;
  logic branch_exec0_is_call_w;
  logic branch_exec0_is_jmp_w;
  logic branch_exec0_is_not_taken_w;
  logic branch_exec0_is_ret_w;
  logic branch_exec0_is_taken_w;
  logic [31:0] branch_exec0_pc_w;
  logic [31:0] branch_exec0_source_w;
  logic branch_exec1_is_call_w;
  logic branch_exec1_is_jmp_w;
  logic branch_exec1_is_not_taken_w;
  logic branch_exec1_is_ret_w;
  logic branch_exec1_is_taken_w;
  logic [31:0] branch_exec1_pc_w;
  logic branch_exec1_request_w;
  logic [31:0] branch_exec1_source_w;
  logic branch_info_is_call_w;
  logic branch_info_is_jmp_w;
  logic branch_info_is_not_taken_w;
  logic branch_info_is_ret_w;
  logic branch_info_is_taken_w;
  logic [31:0] branch_info_pc_w;
  logic branch_info_request_w;
  logic [31:0] branch_info_source_w;
  logic [31:0] branch_pc_w;
  logic branch_request_w;
  input clk_i;
  input [31:0] cpu_id_i;
  logic csr_opcode_invalid_w;
  logic [31:0] csr_opcode_opcode_w;
  logic [31:0] csr_opcode_pc_w;
  logic [4:0] csr_opcode_ra_idx_w;
  logic [31:0] csr_opcode_ra_operand_w;
  logic [4:0] csr_opcode_rb_idx_w;
  logic [31:0] csr_opcode_rb_operand_w;
  logic [4:0] csr_opcode_rd_idx_w;
  logic csr_opcode_valid_w;
  logic [5:0] csr_result_e1_exception_w;
  logic [31:0] csr_result_e1_value_w;
  logic [31:0] csr_result_e1_wdata_w;
  logic csr_result_e1_write_w;
  logic [31:0] csr_writeback_exception_addr_w;
  logic [31:0] csr_writeback_exception_pc_w;
  logic [5:0] csr_writeback_exception_w;
  logic [11:0] csr_writeback_waddr_w;
  logic [31:0] csr_writeback_wdata_w;
  logic csr_writeback_write_w;
  logic div_opcode_valid_w;
  logic exec0_hold_w;
  logic exec0_opcode_valid_w;
  logic exec1_hold_w;
  logic exec1_opcode_valid_w;
  logic fetch0_accept_w;
  logic fetch0_fault_fetch_w;
  logic fetch0_fault_page_w;
  logic fetch0_instr_branch_w;
  logic fetch0_instr_csr_w;
  logic fetch0_instr_div_w;
  logic fetch0_instr_exec_w;
  logic fetch0_instr_invalid_w;
  logic fetch0_instr_lsu_w;
  logic fetch0_instr_mul_w;
  logic fetch0_instr_rd_valid_w;
  logic [31:0] fetch0_instr_w;
  logic [31:0] fetch0_pc_w;
  logic fetch0_valid_w;
  logic fetch1_accept_w;
  logic fetch1_fault_fetch_w;
  logic fetch1_fault_page_w;
  logic fetch1_instr_branch_w;
  logic fetch1_instr_csr_w;
  logic fetch1_instr_div_w;
  logic fetch1_instr_exec_w;
  logic fetch1_instr_invalid_w;
  logic fetch1_instr_lsu_w;
  logic fetch1_instr_mul_w;
  logic fetch1_instr_rd_valid_w;
  logic [31:0] fetch1_instr_w;
  logic [31:0] fetch1_pc_w;
  logic fetch1_valid_w;
  logic ifence_w;
  logic interrupt_inhibit_w;
  input intr_i;
  logic [31:0] lsu_opcode_opcode_w;
  logic [31:0] lsu_opcode_ra_operand_w;
  logic [31:0] lsu_opcode_rb_operand_w;
  logic lsu_opcode_valid_w;
  logic lsu_stall_w;
  input mem_d_accept_i;
  input mem_d_ack_i;
  output [31:0] mem_d_addr_o;
  output mem_d_cacheable_o;
  input [31:0] mem_d_data_rd_i;
  output [31:0] mem_d_data_wr_o;
  input mem_d_error_i;
  output mem_d_flush_o;
  output mem_d_invalidate_o;
  output mem_d_rd_o;
  output [10:0] mem_d_req_tag_o;
  input [10:0] mem_d_resp_tag_i;
  output [3:0] mem_d_wr_o;
  output mem_d_writeback_o;
  input mem_i_accept_i;
  input mem_i_error_i;
  output mem_i_flush_o;
  input [63:0] mem_i_inst_i;
  output mem_i_invalidate_o;
  output [31:0] mem_i_pc_o;
  output mem_i_rd_o;
  input mem_i_valid_i;
  logic mmu_ifetch_accept_w;
  logic mmu_ifetch_error_w;
  logic mmu_ifetch_flush_w;
  logic [63:0] mmu_ifetch_inst_w;
  logic [31:0] mmu_ifetch_pc_w;
  logic mmu_ifetch_rd_w;
  logic mmu_ifetch_valid_w;
  logic mmu_lsu_accept_w;
  logic mmu_lsu_ack_w;
  logic [31:0] mmu_lsu_addr_w;
  logic mmu_lsu_cacheable_w;
  logic [31:0] mmu_lsu_data_rd_w;
  logic [31:0] mmu_lsu_data_wr_w;
  logic mmu_lsu_error_w;
  logic mmu_lsu_flush_w;
  logic mmu_lsu_invalidate_w;
  logic mmu_lsu_rd_w;
  logic [10:0] mmu_lsu_resp_tag_w;
  logic [3:0] mmu_lsu_wr_w;
  logic mmu_lsu_writeback_w;
  logic mmu_mxr_w;
  logic [31:0] mmu_satp_w;
  logic mmu_sum_w;
  logic mul_hold_w;
  logic [31:0] mul_opcode_opcode_w;
  logic [31:0] mul_opcode_ra_operand_w;
  logic [31:0] mul_opcode_rb_operand_w;
  logic mul_opcode_valid_w;
  logic [31:0] opcode0_opcode_w;
  logic [31:0] opcode0_pc_w;
  logic [4:0] opcode0_ra_idx_w;
  logic [31:0] opcode0_ra_operand_w;
  logic [4:0] opcode0_rb_idx_w;
  logic [31:0] opcode0_rb_operand_w;
  logic [4:0] opcode0_rd_idx_w;
  logic [31:0] opcode1_opcode_w;
  logic [31:0] opcode1_pc_w;
  logic [4:0] opcode1_ra_idx_w;
  logic [31:0] opcode1_ra_operand_w;
  logic [4:0] opcode1_rb_idx_w;
  logic [31:0] opcode1_rb_operand_w;
  logic [4:0] opcode1_rd_idx_w;
  input [31:0] reset_vector_i;
  input rst_i;
  logic take_interrupt_w;
  logic [31:0] \u_csr.branch_csr_pc_o ;
  logic \u_csr.branch_csr_request_o ;
  logic \u_csr.branch_q ;
  logic [31:0] \u_csr.branch_target_q ;
  logic \u_csr.clk_i ;
  logic \u_csr.clr_r ;
  logic [31:0] \u_csr.cpu_id_i ;
  logic \u_csr.csr_branch_w ;
  logic [1:0] \u_csr.csr_priv_r ;
  logic [31:0] \u_csr.csr_rdata_w ;
  logic [5:0] \u_csr.csr_result_e1_exception_o ;
  logic [31:0] \u_csr.csr_result_e1_value_o ;
  logic [31:0] \u_csr.csr_result_e1_wdata_o ;
  logic \u_csr.csr_result_e1_write_o ;
  logic [31:0] \u_csr.csr_target_w ;
  logic [31:0] \u_csr.csr_wdata_e1_q ;
  logic \u_csr.csr_write_r ;
  logic [31:0] \u_csr.csr_writeback_exception_addr_i ;
  logic [5:0] \u_csr.csr_writeback_exception_i ;
  logic [31:0] \u_csr.csr_writeback_exception_pc_i ;
  logic [11:0] \u_csr.csr_writeback_waddr_i ;
  logic [31:0] \u_csr.csr_writeback_wdata_i ;
  logic \u_csr.csr_writeback_write_i ;
  logic \u_csr.csrrc_w ;
  logic \u_csr.csrrci_w ;
  logic \u_csr.csrrs_w ;
  logic \u_csr.csrrsi_w ;
  logic \u_csr.csrrw_w ;
  logic \u_csr.csrrwi_w ;
  logic [1:0] \u_csr.current_priv_w ;
  logic [31:0] \u_csr.data_r ;
  logic [5:0] \u_csr.exception_e1_q ;
  logic \u_csr.ifence_o ;
  logic \u_csr.ifence_q ;
  logic \u_csr.ifence_w ;
  logic \u_csr.interrupt_inhibit_i ;
  logic [31:0] \u_csr.interrupt_w ;
  logic \u_csr.intr_i ;
  logic \u_csr.mmu_mxr_o ;
  logic [31:0] \u_csr.mmu_satp_o ;
  logic \u_csr.mmu_sum_o ;
  logic \u_csr.opcode_invalid_i ;
  logic [31:0] \u_csr.opcode_opcode_i ;
  logic [31:0] \u_csr.opcode_pc_i ;
  logic [4:0] \u_csr.opcode_ra_idx_i ;
  logic [31:0] \u_csr.opcode_ra_operand_i ;
  logic [4:0] \u_csr.opcode_rb_idx_i ;
  logic [31:0] \u_csr.opcode_rb_operand_i ;
  logic [4:0] \u_csr.opcode_rd_idx_i ;
  logic \u_csr.opcode_valid_i ;
  logic [31:0] \u_csr.rd_result_e1_q ;
  logic \u_csr.rd_valid_e1_q ;
  logic \u_csr.reset_q ;
  logic [31:0] \u_csr.reset_vector_i ;
  logic \u_csr.rst_i ;
  logic [31:0] \u_csr.satp_reg_w ;
  logic \u_csr.satp_update_w ;
  logic \u_csr.set_r ;
  logic \u_csr.sfence_w ;
  logic [31:0] \u_csr.status_reg_w ;
  logic \u_csr.take_interrupt_o ;
  logic \u_csr.take_interrupt_q ;
  logic \u_csr.u_csrfile.branch_r ;
  logic [31:0] \u_csr.u_csrfile.branch_target_r ;
  logic \u_csr.u_csrfile.buffer_mip_w ;
  logic \u_csr.u_csrfile.clk_i ;
  logic [31:0] \u_csr.u_csrfile.cpu_id_i ;
  logic \u_csr.u_csrfile.csr_branch_o ;
  logic [31:0] \u_csr.u_csrfile.csr_mcause_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mcause_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mcycle_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mcycle_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mepc_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mepc_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mideleg_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mie_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mie_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mip_next_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mip_next_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mip_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mip_r ;
  logic \u_csr.u_csrfile.csr_mip_upd_q ;
  logic [1:0] \u_csr.u_csrfile.csr_mpriv_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mscratch_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mscratch_r ;
  logic \u_csr.u_csrfile.csr_mtime_ie_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mtimecmp_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mtval_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mtval_r ;
  logic [31:0] \u_csr.u_csrfile.csr_mtvec_q ;
  logic [31:0] \u_csr.u_csrfile.csr_mtvec_r ;
  logic [11:0] \u_csr.u_csrfile.csr_raddr_i ;
  logic [31:0] \u_csr.u_csrfile.csr_rdata_o ;
  logic \u_csr.u_csrfile.csr_ren_i ;
  logic [31:0] \u_csr.u_csrfile.csr_satp_q ;
  logic [31:0] \u_csr.u_csrfile.csr_sepc_q ;
  logic [31:0] \u_csr.u_csrfile.csr_sr_q ;
  logic [31:0] \u_csr.u_csrfile.csr_sr_r ;
  logic [31:0] \u_csr.u_csrfile.csr_stvec_q ;
  logic [31:0] \u_csr.u_csrfile.csr_target_o ;
  logic [11:0] \u_csr.u_csrfile.csr_waddr_i ;
  logic [31:0] \u_csr.u_csrfile.csr_wdata_i ;
  logic [31:0] \u_csr.u_csrfile.exception_addr_i ;
  logic [5:0] \u_csr.u_csrfile.exception_i ;
  logic [31:0] \u_csr.u_csrfile.exception_pc_i ;
  logic \u_csr.u_csrfile.ext_intr_i ;
  logic [31:0] \u_csr.u_csrfile.interrupt_o ;
  logic [31:0] \u_csr.u_csrfile.irq_masked_r ;
  logic [31:0] \u_csr.u_csrfile.irq_pending_r ;
  logic [1:0] \u_csr.u_csrfile.irq_priv_q ;
  logic \u_csr.u_csrfile.is_exception_w ;
  logic [1:0] \u_csr.u_csrfile.priv_o ;
  logic [31:0] \u_csr.u_csrfile.rdata_r ;
  logic \u_csr.u_csrfile.rst_i ;
  logic [31:0] \u_csr.u_csrfile.satp_o ;
  logic [31:0] \u_csr.u_csrfile.status_o ;
  logic \u_div.clk_i ;
  logic \u_div.div_busy_q ;
  logic \u_div.div_complete_w ;
  logic \u_div.div_inst_q ;
  logic \u_div.div_operation_w ;
  logic \u_div.div_rem_inst_w ;
  logic [31:0] \u_div.div_result_r ;
  logic \u_div.div_start_w ;
  logic [31:0] \u_div.dividend_q ;
  logic [62:0] \u_div.divisor_q ;
  logic \u_div.inst_div_w ;
  logic \u_div.inst_divu_w ;
  logic \u_div.inst_rem_w ;
  logic \u_div.inst_remu_w ;
  logic \u_div.invert_res_q ;
  logic [31:0] \u_div.last_a_q ;
  logic [31:0] \u_div.last_b_q ;
  logic \u_div.last_div_q ;
  logic \u_div.last_divu_q ;
  logic \u_div.last_rem_q ;
  logic \u_div.last_remu_q ;
  logic [31:0] \u_div.opcode_opcode_i ;
  logic [31:0] \u_div.opcode_pc_i ;
  logic [4:0] \u_div.opcode_ra_idx_i ;
  logic [31:0] \u_div.opcode_ra_operand_i ;
  logic [4:0] \u_div.opcode_rb_idx_i ;
  logic [31:0] \u_div.opcode_rb_operand_i ;
  logic [4:0] \u_div.opcode_rd_idx_i ;
  logic \u_div.opcode_valid_i ;
  logic [31:0] \u_div.q_mask_q ;
  logic [31:0] \u_div.quotient_q ;
  logic \u_div.rst_i ;
  logic \u_div.signed_operation_w ;
  logic \u_div.valid_q ;
  logic [31:0] \u_div.wb_result_q ;
  logic \u_div.writeback_valid_o ;
  logic [31:0] \u_div.writeback_value_o ;
  logic [3:0] \u_exec0.alu_func_r ;
  logic [31:0] \u_exec0.alu_input_a_r ;
  logic [31:0] \u_exec0.alu_input_b_r ;
  logic [31:0] \u_exec0.alu_p_w ;
  logic [31:0] \u_exec0.bimm_r ;
  logic \u_exec0.branch_call_q ;
  logic \u_exec0.branch_call_r ;
  logic [31:0] \u_exec0.branch_d_pc_o ;
  logic \u_exec0.branch_d_request_o ;
  logic \u_exec0.branch_is_call_o ;
  logic \u_exec0.branch_is_jmp_o ;
  logic \u_exec0.branch_is_not_taken_o ;
  logic \u_exec0.branch_is_ret_o ;
  logic \u_exec0.branch_is_taken_o ;
  logic \u_exec0.branch_jmp_q ;
  logic \u_exec0.branch_jmp_r ;
  logic \u_exec0.branch_ntaken_q ;
  logic [31:0] \u_exec0.branch_pc_o ;
  logic \u_exec0.branch_r ;
  logic \u_exec0.branch_ret_q ;
  logic \u_exec0.branch_ret_r ;
  logic [31:0] \u_exec0.branch_source_o ;
  logic \u_exec0.branch_taken_q ;
  logic \u_exec0.branch_taken_r ;
  logic [31:0] \u_exec0.branch_target_r ;
  logic \u_exec0.clk_i ;
  logic \u_exec0.hold_i ;
  logic [31:0] \u_exec0.imm12_r ;
  logic [31:0] \u_exec0.imm20_r ;
  logic [31:0] \u_exec0.jimm20_r ;
  logic [31:0] \u_exec0.opcode_opcode_i ;
  logic [31:0] \u_exec0.opcode_pc_i ;
  logic [4:0] \u_exec0.opcode_ra_idx_i ;
  logic [31:0] \u_exec0.opcode_ra_operand_i ;
  logic [4:0] \u_exec0.opcode_rb_idx_i ;
  logic [31:0] \u_exec0.opcode_rb_operand_i ;
  logic [4:0] \u_exec0.opcode_rd_idx_i ;
  logic \u_exec0.opcode_valid_i ;
  logic [31:0] \u_exec0.pc_m_q ;
  logic [31:0] \u_exec0.pc_x_q ;
  logic [31:0] \u_exec0.result_q ;
  logic \u_exec0.rst_i ;
  logic [4:0] \u_exec0.shamt_r ;
  logic [31:0] \u_exec0.u_alu.alu_a_i ;
  logic [31:0] \u_exec0.u_alu.alu_b_i ;
  logic [3:0] \u_exec0.u_alu.alu_op_i ;
  logic [31:0] \u_exec0.u_alu.alu_p_o ;
  logic [31:0] \u_exec0.u_alu.result_r ;
  logic [31:0] \u_exec0.u_alu.sub_res_w ;
  logic [31:0] \u_exec0.writeback_value_o ;
  logic [3:0] \u_exec1.alu_func_r ;
  logic [31:0] \u_exec1.alu_input_a_r ;
  logic [31:0] \u_exec1.alu_input_b_r ;
  logic [31:0] \u_exec1.alu_p_w ;
  logic [31:0] \u_exec1.bimm_r ;
  logic \u_exec1.branch_call_q ;
  logic \u_exec1.branch_call_r ;
  logic [31:0] \u_exec1.branch_d_pc_o ;
  logic \u_exec1.branch_d_request_o ;
  logic \u_exec1.branch_is_call_o ;
  logic \u_exec1.branch_is_jmp_o ;
  logic \u_exec1.branch_is_not_taken_o ;
  logic \u_exec1.branch_is_ret_o ;
  logic \u_exec1.branch_is_taken_o ;
  logic \u_exec1.branch_jmp_q ;
  logic \u_exec1.branch_jmp_r ;
  logic \u_exec1.branch_ntaken_q ;
  logic [31:0] \u_exec1.branch_pc_o ;
  logic \u_exec1.branch_r ;
  logic \u_exec1.branch_request_o ;
  logic \u_exec1.branch_ret_q ;
  logic \u_exec1.branch_ret_r ;
  logic [31:0] \u_exec1.branch_source_o ;
  logic \u_exec1.branch_taken_q ;
  logic \u_exec1.branch_taken_r ;
  logic [31:0] \u_exec1.branch_target_r ;
  logic \u_exec1.clk_i ;
  logic \u_exec1.hold_i ;
  logic [31:0] \u_exec1.imm12_r ;
  logic [31:0] \u_exec1.imm20_r ;
  logic [31:0] \u_exec1.jimm20_r ;
  logic [31:0] \u_exec1.opcode_opcode_i ;
  logic [31:0] \u_exec1.opcode_pc_i ;
  logic [4:0] \u_exec1.opcode_ra_idx_i ;
  logic [31:0] \u_exec1.opcode_ra_operand_i ;
  logic [4:0] \u_exec1.opcode_rb_idx_i ;
  logic [31:0] \u_exec1.opcode_rb_operand_i ;
  logic [4:0] \u_exec1.opcode_rd_idx_i ;
  logic \u_exec1.opcode_valid_i ;
  logic [31:0] \u_exec1.pc_m_q ;
  logic [31:0] \u_exec1.pc_x_q ;
  logic [31:0] \u_exec1.result_q ;
  logic \u_exec1.rst_i ;
  logic [4:0] \u_exec1.shamt_r ;
  logic [31:0] \u_exec1.u_alu.alu_a_i ;
  logic [31:0] \u_exec1.u_alu.alu_b_i ;
  logic [3:0] \u_exec1.u_alu.alu_op_i ;
  logic [31:0] \u_exec1.u_alu.alu_p_o ;
  logic [31:0] \u_exec1.u_alu.result_r ;
  logic [31:0] \u_exec1.u_alu.sub_res_w ;
  logic [31:0] \u_exec1.writeback_value_o ;
  logic \u_frontend.branch_info_is_call_i ;
  logic \u_frontend.branch_info_is_jmp_i ;
  logic \u_frontend.branch_info_is_not_taken_i ;
  logic \u_frontend.branch_info_is_ret_i ;
  logic \u_frontend.branch_info_is_taken_i ;
  logic [31:0] \u_frontend.branch_info_pc_i ;
  logic \u_frontend.branch_info_request_i ;
  logic [31:0] \u_frontend.branch_info_source_i ;
  logic [31:0] \u_frontend.branch_pc_i ;
  logic \u_frontend.branch_request_i ;
  logic \u_frontend.clk_i ;
  logic \u_frontend.fetch0_accept_i ;
  logic \u_frontend.fetch0_fault_fetch_o ;
  logic \u_frontend.fetch0_fault_page_o ;
  logic \u_frontend.fetch0_instr_branch_o ;
  logic \u_frontend.fetch0_instr_csr_o ;
  logic \u_frontend.fetch0_instr_div_o ;
  logic \u_frontend.fetch0_instr_exec_o ;
  logic \u_frontend.fetch0_instr_invalid_o ;
  logic \u_frontend.fetch0_instr_lsu_o ;
  logic \u_frontend.fetch0_instr_mul_o ;
  logic [31:0] \u_frontend.fetch0_instr_o ;
  logic \u_frontend.fetch0_instr_rd_valid_o ;
  logic [31:0] \u_frontend.fetch0_pc_o ;
  logic \u_frontend.fetch0_valid_o ;
  logic \u_frontend.fetch1_accept_i ;
  logic \u_frontend.fetch1_fault_fetch_o ;
  logic \u_frontend.fetch1_fault_page_o ;
  logic \u_frontend.fetch1_instr_branch_o ;
  logic \u_frontend.fetch1_instr_csr_o ;
  logic \u_frontend.fetch1_instr_div_o ;
  logic \u_frontend.fetch1_instr_exec_o ;
  logic \u_frontend.fetch1_instr_invalid_o ;
  logic \u_frontend.fetch1_instr_lsu_o ;
  logic \u_frontend.fetch1_instr_mul_o ;
  logic [31:0] \u_frontend.fetch1_instr_o ;
  logic \u_frontend.fetch1_instr_rd_valid_o ;
  logic [31:0] \u_frontend.fetch1_pc_o ;
  logic \u_frontend.fetch1_valid_o ;
  logic \u_frontend.fetch_accept_w ;
  logic \u_frontend.fetch_fault_fetch_w ;
  logic \u_frontend.fetch_fault_page_w ;
  logic [63:0] \u_frontend.fetch_instr_w ;
  logic \u_frontend.fetch_invalidate_i ;
  logic \u_frontend.fetch_pc_accept_w ;
  logic [31:0] \u_frontend.fetch_pc_f_w ;
  logic [31:0] \u_frontend.fetch_pc_w ;
  logic [1:0] \u_frontend.fetch_pred_branch_w ;
  logic \u_frontend.fetch_valid_w ;
  logic \u_frontend.icache_accept_i ;
  logic \u_frontend.icache_error_i ;
  logic \u_frontend.icache_flush_o ;
  logic [63:0] \u_frontend.icache_inst_i ;
  logic [31:0] \u_frontend.icache_pc_o ;
  logic \u_frontend.icache_rd_o ;
  logic \u_frontend.icache_valid_i ;
  logic [31:0] \u_frontend.next_pc_f_w ;
  logic [1:0] \u_frontend.next_taken_f_w ;
  logic \u_frontend.rst_i ;
  logic [31:0] \u_frontend.u_decode.branch_pc_i ;
  logic \u_frontend.u_decode.branch_request_i ;
  logic \u_frontend.u_decode.clk_i ;
  logic \u_frontend.u_decode.fetch_in_accept_o ;
  logic \u_frontend.u_decode.fetch_in_fault_fetch_i ;
  logic \u_frontend.u_decode.fetch_in_fault_page_i ;
  logic [63:0] \u_frontend.u_decode.fetch_in_instr_i ;
  logic [31:0] \u_frontend.u_decode.fetch_in_pc_i ;
  logic [1:0] \u_frontend.u_decode.fetch_in_pred_branch_i ;
  logic \u_frontend.u_decode.fetch_in_valid_i ;
  logic \u_frontend.u_decode.fetch_out0_accept_i ;
  logic \u_frontend.u_decode.fetch_out0_fault_fetch_o ;
  logic \u_frontend.u_decode.fetch_out0_fault_page_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_branch_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_csr_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_div_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_exec_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_invalid_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_lsu_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_mul_o ;
  logic [31:0] \u_frontend.u_decode.fetch_out0_instr_o ;
  logic \u_frontend.u_decode.fetch_out0_instr_rd_valid_o ;
  logic [31:0] \u_frontend.u_decode.fetch_out0_pc_o ;
  logic \u_frontend.u_decode.fetch_out0_valid_o ;
  logic \u_frontend.u_decode.fetch_out1_accept_i ;
  logic \u_frontend.u_decode.fetch_out1_fault_fetch_o ;
  logic \u_frontend.u_decode.fetch_out1_fault_page_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_branch_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_csr_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_div_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_exec_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_invalid_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_lsu_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_mul_o ;
  logic [31:0] \u_frontend.u_decode.fetch_out1_instr_o ;
  logic \u_frontend.u_decode.fetch_out1_instr_rd_valid_o ;
  logic [31:0] \u_frontend.u_decode.fetch_out1_pc_o ;
  logic \u_frontend.u_decode.fetch_out1_valid_o ;
  logic \u_frontend.u_decode.rst_i ;
  logic \u_frontend.u_decode.u_dec0.branch_o ;
  logic \u_frontend.u_decode.u_dec0.csr_o ;
  logic \u_frontend.u_decode.u_dec0.div_o ;
  logic \u_frontend.u_decode.u_dec0.exec_o ;
  logic \u_frontend.u_decode.u_dec0.fetch_fault_i ;
  logic \u_frontend.u_decode.u_dec0.invalid_o ;
  logic \u_frontend.u_decode.u_dec0.invalid_w ;
  logic \u_frontend.u_decode.u_dec0.lsu_o ;
  logic \u_frontend.u_decode.u_dec0.mul_o ;
  logic [31:0] \u_frontend.u_decode.u_dec0.opcode_i ;
  logic \u_frontend.u_decode.u_dec0.rd_valid_o ;
  logic \u_frontend.u_decode.u_dec0.valid_i ;
  logic \u_frontend.u_decode.u_dec1.branch_o ;
  logic \u_frontend.u_decode.u_dec1.csr_o ;
  logic \u_frontend.u_decode.u_dec1.div_o ;
  logic \u_frontend.u_decode.u_dec1.exec_o ;
  logic \u_frontend.u_decode.u_dec1.fetch_fault_i ;
  logic \u_frontend.u_decode.u_dec1.invalid_o ;
  logic \u_frontend.u_decode.u_dec1.invalid_w ;
  logic \u_frontend.u_decode.u_dec1.lsu_o ;
  logic \u_frontend.u_decode.u_dec1.mul_o ;
  logic [31:0] \u_frontend.u_decode.u_dec1.opcode_i ;
  logic \u_frontend.u_decode.u_dec1.rd_valid_o ;
  logic \u_frontend.u_decode.u_dec1.valid_i ;
  logic \u_frontend.u_decode.u_fifo.accept_o ;
  logic \u_frontend.u_decode.u_fifo.clk_i ;
  logic [1:0] \u_frontend.u_decode.u_fifo.count_q ;
  logic [31:0] \u_frontend.u_decode.u_fifo.data0_out_o ;
  logic [31:0] \u_frontend.u_decode.u_fifo.data1_out_o ;
  logic [63:0] \u_frontend.u_decode.u_fifo.data_in_i ;
  logic \u_frontend.u_decode.u_fifo.flush_i ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info0_in_i ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info0_out_o ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info0_q[0] ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info0_q[1] ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info1_in_i ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info1_out_o ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info1_q[0] ;
  logic [1:0] \u_frontend.u_decode.u_fifo.info1_q[1] ;
  logic [31:0] \u_frontend.u_decode.u_fifo.pc0_out_o ;
  logic [31:0] \u_frontend.u_decode.u_fifo.pc1_out_o ;
  logic [31:0] \u_frontend.u_decode.u_fifo.pc_in_i ;
  logic [31:0] \u_frontend.u_decode.u_fifo.pc_q[0] ;
  logic [31:0] \u_frontend.u_decode.u_fifo.pc_q[1] ;
  logic \u_frontend.u_decode.u_fifo.pop0_i ;
  logic \u_frontend.u_decode.u_fifo.pop1_i ;
  logic \u_frontend.u_decode.u_fifo.pop1_w ;
  logic \u_frontend.u_decode.u_fifo.pop2_w ;
  logic \u_frontend.u_decode.u_fifo.pop_complete_w ;
  logic [1:0] \u_frontend.u_decode.u_fifo.pred_in_i ;
  logic \u_frontend.u_decode.u_fifo.push_i ;
  logic \u_frontend.u_decode.u_fifo.push_w ;
  logic [63:0] \u_frontend.u_decode.u_fifo.ram_q[0] ;
  logic [63:0] \u_frontend.u_decode.u_fifo.ram_q[1] ;
  logic \u_frontend.u_decode.u_fifo.rd_ptr_q ;
  logic \u_frontend.u_decode.u_fifo.rst_i ;
  logic \u_frontend.u_decode.u_fifo.valid0_o ;
  logic \u_frontend.u_decode.u_fifo.valid0_q[0] ;
  logic \u_frontend.u_decode.u_fifo.valid0_q[1] ;
  logic \u_frontend.u_decode.u_fifo.valid1_o ;
  logic \u_frontend.u_decode.u_fifo.valid1_q[0] ;
  logic \u_frontend.u_decode.u_fifo.valid1_q[1] ;
  logic \u_frontend.u_decode.u_fifo.wr_ptr_q ;
  logic \u_frontend.u_fetch.active_q ;
  logic [31:0] \u_frontend.u_fetch.branch_pc_i ;
  logic [31:0] \u_frontend.u_fetch.branch_pc_q ;
  logic [31:0] \u_frontend.u_fetch.branch_pc_w ;
  logic \u_frontend.u_fetch.branch_q ;
  logic \u_frontend.u_fetch.branch_request_i ;
  logic \u_frontend.u_fetch.branch_w ;
  logic \u_frontend.u_fetch.clk_i ;
  logic \u_frontend.u_fetch.fetch_accept_i ;
  logic \u_frontend.u_fetch.fetch_fault_fetch_o ;
  logic \u_frontend.u_fetch.fetch_fault_page_o ;
  logic [63:0] \u_frontend.u_fetch.fetch_instr_o ;
  logic \u_frontend.u_fetch.fetch_invalidate_i ;
  logic [31:0] \u_frontend.u_fetch.fetch_pc_o ;
  logic [1:0] \u_frontend.u_fetch.fetch_pred_branch_o ;
  logic \u_frontend.u_fetch.fetch_resp_drop_w ;
  logic \u_frontend.u_fetch.fetch_valid_o ;
  logic \u_frontend.u_fetch.icache_accept_i ;
  logic \u_frontend.u_fetch.icache_busy_w ;
  logic \u_frontend.u_fetch.icache_error_i ;
  logic \u_frontend.u_fetch.icache_fetch_q ;
  logic \u_frontend.u_fetch.icache_flush_o ;
  logic [63:0] \u_frontend.u_fetch.icache_inst_i ;
  logic \u_frontend.u_fetch.icache_invalidate_q ;
  logic [31:0] \u_frontend.u_fetch.icache_pc_o ;
  logic [31:0] \u_frontend.u_fetch.icache_pc_w ;
  logic \u_frontend.u_fetch.icache_rd_o ;
  logic \u_frontend.u_fetch.icache_valid_i ;
  logic [31:0] \u_frontend.u_fetch.next_pc_f_i ;
  logic [1:0] \u_frontend.u_fetch.next_taken_f_i ;
  logic \u_frontend.u_fetch.pc_accept_o ;
  logic [31:0] \u_frontend.u_fetch.pc_d_q ;
  logic [31:0] \u_frontend.u_fetch.pc_f_o ;
  logic [31:0] \u_frontend.u_fetch.pc_f_q ;
  logic [1:0] \u_frontend.u_fetch.pred_d_q ;
  logic \u_frontend.u_fetch.rst_i ;
  logic [99:0] \u_frontend.u_fetch.skid_buffer_q ;
  logic \u_frontend.u_fetch.skid_valid_q ;
  logic \u_frontend.u_fetch.stall_q ;
  logic \u_frontend.u_fetch.stall_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.bht_predict_taken_w ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_rd_entry_w ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[0] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[1] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[2] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[3] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[4] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[5] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[6] ;
  logic [1:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[7] ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.bht_wr_entry_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_hit_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_miss_r ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_next_pc_r ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_w ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_alloc_w ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.ras_call_pred_w ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_q ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_r ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_pc_pred_w ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.ras_ret_pred_w ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[0] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[1] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[2] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[3] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[4] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[5] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[6] ;
  logic [31:0] \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[7] ;
  logic [2:0] \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.alloc_entry_o ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.alloc_i ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.clk_i ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.hit_i ;
  logic [15:0] \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q ;
  logic \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.rst_i ;
  logic \u_frontend.u_npc.branch_is_call_i ;
  logic \u_frontend.u_npc.branch_is_jmp_i ;
  logic \u_frontend.u_npc.branch_is_not_taken_i ;
  logic \u_frontend.u_npc.branch_is_ret_i ;
  logic \u_frontend.u_npc.branch_is_taken_i ;
  logic [31:0] \u_frontend.u_npc.branch_pc_i ;
  logic \u_frontend.u_npc.branch_request_i ;
  logic [31:0] \u_frontend.u_npc.branch_source_i ;
  logic \u_frontend.u_npc.clk_i ;
  logic [31:0] \u_frontend.u_npc.next_pc_f_o ;
  logic [1:0] \u_frontend.u_npc.next_taken_f_o ;
  logic \u_frontend.u_npc.pc_accept_i ;
  logic [31:0] \u_frontend.u_npc.pc_f_i ;
  logic \u_frontend.u_npc.rst_i ;
  logic [31:0] \u_issue.branch_csr_pc_i ;
  logic \u_issue.branch_csr_request_i ;
  logic [31:0] \u_issue.branch_d_exec0_pc_i ;
  logic \u_issue.branch_d_exec0_request_i ;
  logic [31:0] \u_issue.branch_d_exec1_pc_i ;
  logic \u_issue.branch_d_exec1_request_i ;
  logic \u_issue.branch_exec0_is_call_i ;
  logic \u_issue.branch_exec0_is_jmp_i ;
  logic \u_issue.branch_exec0_is_not_taken_i ;
  logic \u_issue.branch_exec0_is_ret_i ;
  logic \u_issue.branch_exec0_is_taken_i ;
  logic [31:0] \u_issue.branch_exec0_pc_i ;
  logic [31:0] \u_issue.branch_exec0_source_i ;
  logic \u_issue.branch_exec1_is_call_i ;
  logic \u_issue.branch_exec1_is_jmp_i ;
  logic \u_issue.branch_exec1_is_not_taken_i ;
  logic \u_issue.branch_exec1_is_ret_i ;
  logic \u_issue.branch_exec1_is_taken_i ;
  logic [31:0] \u_issue.branch_exec1_pc_i ;
  logic \u_issue.branch_exec1_request_i ;
  logic [31:0] \u_issue.branch_exec1_source_i ;
  logic \u_issue.branch_info_is_call_o ;
  logic \u_issue.branch_info_is_jmp_o ;
  logic \u_issue.branch_info_is_not_taken_o ;
  logic \u_issue.branch_info_is_ret_o ;
  logic \u_issue.branch_info_is_taken_o ;
  logic [31:0] \u_issue.branch_info_pc_o ;
  logic \u_issue.branch_info_request_o ;
  logic [31:0] \u_issue.branch_info_source_o ;
  logic [31:0] \u_issue.branch_pc_o ;
  logic \u_issue.branch_request_o ;
  logic \u_issue.clk_i ;
  logic \u_issue.csr_opcode_invalid_o ;
  logic [31:0] \u_issue.csr_opcode_opcode_o ;
  logic [31:0] \u_issue.csr_opcode_pc_o ;
  logic [4:0] \u_issue.csr_opcode_ra_idx_o ;
  logic [31:0] \u_issue.csr_opcode_ra_operand_o ;
  logic [4:0] \u_issue.csr_opcode_rb_idx_o ;
  logic [31:0] \u_issue.csr_opcode_rb_operand_o ;
  logic [4:0] \u_issue.csr_opcode_rd_idx_o ;
  logic \u_issue.csr_opcode_valid_o ;
  logic \u_issue.csr_pending_q ;
  logic [5:0] \u_issue.csr_result_e1_exception_i ;
  logic [31:0] \u_issue.csr_result_e1_value_i ;
  logic [31:0] \u_issue.csr_result_e1_wdata_i ;
  logic \u_issue.csr_result_e1_write_i ;
  logic [31:0] \u_issue.csr_writeback_exception_addr_o ;
  logic [5:0] \u_issue.csr_writeback_exception_o ;
  logic [31:0] \u_issue.csr_writeback_exception_pc_o ;
  logic [11:0] \u_issue.csr_writeback_waddr_o ;
  logic [31:0] \u_issue.csr_writeback_wdata_o ;
  logic \u_issue.csr_writeback_write_o ;
  logic \u_issue.div_opcode_valid_o ;
  logic \u_issue.div_pending_q ;
  logic \u_issue.dual_issue_ok_w ;
  logic \u_issue.dual_issue_w ;
  logic \u_issue.exec0_hold_o ;
  logic \u_issue.exec0_opcode_valid_o ;
  logic \u_issue.exec1_hold_o ;
  logic \u_issue.exec1_opcode_valid_o ;
  logic \u_issue.fetch0_accept_o ;
  logic \u_issue.fetch0_fault_fetch_i ;
  logic \u_issue.fetch0_fault_page_i ;
  logic \u_issue.fetch0_instr_branch_i ;
  logic \u_issue.fetch0_instr_csr_i ;
  logic \u_issue.fetch0_instr_div_i ;
  logic \u_issue.fetch0_instr_exec_i ;
  logic [31:0] \u_issue.fetch0_instr_i ;
  logic \u_issue.fetch0_instr_invalid_i ;
  logic \u_issue.fetch0_instr_lsu_i ;
  logic \u_issue.fetch0_instr_mul_i ;
  logic \u_issue.fetch0_instr_rd_valid_i ;
  logic [31:0] \u_issue.fetch0_pc_i ;
  logic \u_issue.fetch0_valid_i ;
  logic \u_issue.fetch1_accept_o ;
  logic \u_issue.fetch1_fault_fetch_i ;
  logic \u_issue.fetch1_fault_page_i ;
  logic \u_issue.fetch1_instr_branch_i ;
  logic \u_issue.fetch1_instr_csr_i ;
  logic \u_issue.fetch1_instr_div_i ;
  logic \u_issue.fetch1_instr_exec_i ;
  logic [31:0] \u_issue.fetch1_instr_i ;
  logic \u_issue.fetch1_instr_invalid_i ;
  logic \u_issue.fetch1_instr_lsu_i ;
  logic \u_issue.fetch1_instr_mul_i ;
  logic \u_issue.fetch1_instr_rd_valid_i ;
  logic [31:0] \u_issue.fetch1_pc_i ;
  logic \u_issue.fetch1_valid_i ;
  logic \u_issue.interrupt_inhibit_o ;
  logic \u_issue.issue_a_branch_w ;
  logic \u_issue.issue_a_csr_w ;
  logic \u_issue.issue_a_div_w ;
  logic \u_issue.issue_a_exec_w ;
  logic [4:0] \u_issue.issue_a_fault_w ;
  logic \u_issue.issue_a_invalid_w ;
  logic \u_issue.issue_a_lsu_w ;
  logic \u_issue.issue_a_mul_w ;
  logic [4:0] \u_issue.issue_a_ra_idx_w ;
  logic [31:0] \u_issue.issue_a_ra_value_r ;
  logic [31:0] \u_issue.issue_a_ra_value_w ;
  logic [4:0] \u_issue.issue_a_rb_idx_w ;
  logic [31:0] \u_issue.issue_a_rb_value_r ;
  logic [31:0] \u_issue.issue_a_rb_value_w ;
  logic [4:0] \u_issue.issue_a_rd_idx_w ;
  logic \u_issue.issue_a_sb_alloc_w ;
  logic \u_issue.issue_b_branch_w ;
  logic \u_issue.issue_b_csr_w ;
  logic \u_issue.issue_b_div_w ;
  logic \u_issue.issue_b_exec_w ;
  logic [4:0] \u_issue.issue_b_fault_w ;
  logic \u_issue.issue_b_invalid_w ;
  logic \u_issue.issue_b_lsu_w ;
  logic \u_issue.issue_b_mul_w ;
  logic [4:0] \u_issue.issue_b_ra_idx_w ;
  logic [31:0] \u_issue.issue_b_ra_value_r ;
  logic [31:0] \u_issue.issue_b_ra_value_w ;
  logic [4:0] \u_issue.issue_b_rb_idx_w ;
  logic [31:0] \u_issue.issue_b_rb_value_r ;
  logic [31:0] \u_issue.issue_b_rb_value_w ;
  logic [4:0] \u_issue.issue_b_rd_idx_w ;
  logic \u_issue.issue_b_sb_alloc_w ;
  logic [31:0] \u_issue.lsu_opcode_opcode_o ;
  logic [31:0] \u_issue.lsu_opcode_ra_operand_o ;
  logic [31:0] \u_issue.lsu_opcode_rb_operand_o ;
  logic \u_issue.lsu_opcode_valid_o ;
  logic \u_issue.lsu_stall_i ;
  logic \u_issue.mispredicted_r ;
  logic \u_issue.mul_hold_o ;
  logic [31:0] \u_issue.mul_opcode_opcode_o ;
  logic [31:0] \u_issue.mul_opcode_ra_operand_o ;
  logic [31:0] \u_issue.mul_opcode_rb_operand_o ;
  logic \u_issue.mul_opcode_valid_o ;
  logic [31:0] \u_issue.opcode0_opcode_o ;
  logic [31:0] \u_issue.opcode0_pc_o ;
  logic [4:0] \u_issue.opcode0_ra_idx_o ;
  logic [31:0] \u_issue.opcode0_ra_operand_o ;
  logic [4:0] \u_issue.opcode0_rb_idx_o ;
  logic [31:0] \u_issue.opcode0_rb_operand_o ;
  logic [4:0] \u_issue.opcode0_rd_idx_o ;
  logic [31:0] \u_issue.opcode1_opcode_o ;
  logic [31:0] \u_issue.opcode1_pc_o ;
  logic [4:0] \u_issue.opcode1_ra_idx_o ;
  logic [31:0] \u_issue.opcode1_ra_operand_o ;
  logic [4:0] \u_issue.opcode1_rb_idx_o ;
  logic [31:0] \u_issue.opcode1_rb_operand_o ;
  logic [4:0] \u_issue.opcode1_rd_idx_o ;
  logic \u_issue.opcode_a_accept_r ;
  logic [1:0] \u_issue.opcode_a_fault_r ;
  logic \u_issue.opcode_a_issue_r ;
  logic [31:0] \u_issue.opcode_a_pc_r ;
  logic [31:0] \u_issue.opcode_a_r ;
  logic \u_issue.opcode_a_valid_r ;
  logic \u_issue.opcode_b_accept_r ;
  logic [1:0] \u_issue.opcode_b_fault_r ;
  logic \u_issue.opcode_b_issue_r ;
  logic [31:0] \u_issue.opcode_b_pc_r ;
  logic [31:0] \u_issue.opcode_b_r ;
  logic \u_issue.opcode_b_valid_r ;
  logic [31:0] \u_issue.pc_x_q ;
  logic \u_issue.pipe0_branch_e1_w ;
  logic \u_issue.pipe0_csr_wb_w ;
  logic [5:0] \u_issue.pipe0_exception_wb_w ;
  logic \u_issue.pipe0_load_e1_w ;
  logic \u_issue.pipe0_load_e2_w ;
  logic \u_issue.pipe0_mul_e1_w ;
  logic \u_issue.pipe0_mul_e2_w ;
  logic [31:0] \u_issue.pipe0_opc_wb_w ;
  logic [31:0] \u_issue.pipe0_opcode_e1_w ;
  logic [31:0] \u_issue.pipe0_pc_e1_w ;
  logic [31:0] \u_issue.pipe0_pc_wb_w ;
  logic [4:0] \u_issue.pipe0_rd_e1_w ;
  logic [4:0] \u_issue.pipe0_rd_e2_w ;
  logic [4:0] \u_issue.pipe0_rd_wb_w ;
  logic [31:0] \u_issue.pipe0_result_e2_w ;
  logic [31:0] \u_issue.pipe0_result_wb_w ;
  logic \u_issue.pipe0_squash_e1_e2_w ;
  logic \u_issue.pipe0_stall_raw_w ;
  logic \u_issue.pipe0_store_e1_w ;
  logic \u_issue.pipe0_valid_wb_w ;
  logic \u_issue.pipe1_branch_e1_w ;
  logic [5:0] \u_issue.pipe1_exception_wb_w ;
  logic \u_issue.pipe1_load_e1_w ;
  logic \u_issue.pipe1_load_e2_w ;
  logic \u_issue.pipe1_mul_e1_w ;
  logic \u_issue.pipe1_mul_e2_w ;
  logic \u_issue.pipe1_mux_lsu_r ;
  logic \u_issue.pipe1_mux_mul_r ;
  logic \u_issue.pipe1_ok_w ;
  logic [31:0] \u_issue.pipe1_opc_wb_w ;
  logic [31:0] \u_issue.pipe1_opcode_e1_w ;
  logic [31:0] \u_issue.pipe1_pc_e1_w ;
  logic [31:0] \u_issue.pipe1_pc_wb_w ;
  logic [4:0] \u_issue.pipe1_rd_e1_w ;
  logic [4:0] \u_issue.pipe1_rd_e2_w ;
  logic [4:0] \u_issue.pipe1_rd_wb_w ;
  logic [31:0] \u_issue.pipe1_result_e2_w ;
  logic [31:0] \u_issue.pipe1_result_wb_w ;
  logic \u_issue.pipe1_squash_e1_e2_w ;
  logic \u_issue.pipe1_stall_raw_w ;
  logic \u_issue.pipe1_store_e1_w ;
  logic \u_issue.pipe1_valid_wb_w ;
  logic \u_issue.rst_i ;
  logic \u_issue.single_issue_w ;
  logic \u_issue.slot0_valid_r ;
  logic \u_issue.slot1_valid_r ;
  logic \u_issue.squash_w ;
  logic \u_issue.stall_w ;
  logic \u_issue.take_interrupt_i ;
  logic \u_issue.u_pipe0_ctrl.alu_e1_w ;
  logic [31:0] \u_issue.u_pipe0_ctrl.alu_result_e1_i ;
  logic \u_issue.u_pipe0_ctrl.branch_e1_o ;
  logic \u_issue.u_pipe0_ctrl.branch_misaligned_w ;
  logic \u_issue.u_pipe0_ctrl.clk_i ;
  logic \u_issue.u_pipe0_ctrl.csr_e1_w ;
  logic [5:0] \u_issue.u_pipe0_ctrl.csr_result_exception_e1_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.csr_result_value_e1_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.csr_result_wdata_e1_i ;
  logic \u_issue.u_pipe0_ctrl.csr_result_write_e1_i ;
  logic [11:0] \u_issue.u_pipe0_ctrl.csr_waddr_wb_o ;
  logic \u_issue.u_pipe0_ctrl.csr_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.csr_wdata_e2_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.csr_wdata_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  logic \u_issue.u_pipe0_ctrl.csr_wr_e2_q ;
  logic \u_issue.u_pipe0_ctrl.csr_wr_wb_q ;
  logic \u_issue.u_pipe0_ctrl.csr_write_wb_o ;
  logic [9:0] \u_issue.u_pipe0_ctrl.ctrl_e1_q ;
  logic [9:0] \u_issue.u_pipe0_ctrl.ctrl_e2_q ;
  logic [9:0] \u_issue.u_pipe0_ctrl.ctrl_wb_q ;
  logic \u_issue.u_pipe0_ctrl.div_complete_i ;
  logic \u_issue.u_pipe0_ctrl.div_e1_w ;
  logic [31:0] \u_issue.u_pipe0_ctrl.div_result_i ;
  logic [5:0] \u_issue.u_pipe0_ctrl.exception_e1_q ;
  logic [5:0] \u_issue.u_pipe0_ctrl.exception_e2_q ;
  logic [5:0] \u_issue.u_pipe0_ctrl.exception_e2_r ;
  logic [5:0] \u_issue.u_pipe0_ctrl.exception_wb_o ;
  logic [5:0] \u_issue.u_pipe0_ctrl.exception_wb_q ;
  logic \u_issue.u_pipe0_ctrl.issue_accept_i ;
  logic \u_issue.u_pipe0_ctrl.issue_branch_i ;
  logic \u_issue.u_pipe0_ctrl.issue_branch_taken_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.issue_branch_target_i ;
  logic \u_issue.u_pipe0_ctrl.issue_csr_i ;
  logic \u_issue.u_pipe0_ctrl.issue_div_i ;
  logic [5:0] \u_issue.u_pipe0_ctrl.issue_exception_i ;
  logic \u_issue.u_pipe0_ctrl.issue_lsu_i ;
  logic \u_issue.u_pipe0_ctrl.issue_mul_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.issue_opcode_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.issue_operand_ra_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.issue_operand_rb_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.issue_pc_i ;
  logic [4:0] \u_issue.u_pipe0_ctrl.issue_rd_i ;
  logic \u_issue.u_pipe0_ctrl.issue_rd_valid_i ;
  logic \u_issue.u_pipe0_ctrl.issue_stall_i ;
  logic \u_issue.u_pipe0_ctrl.issue_valid_i ;
  logic \u_issue.u_pipe0_ctrl.load_e1_o ;
  logic \u_issue.u_pipe0_ctrl.load_e2_o ;
  logic \u_issue.u_pipe0_ctrl.mem_complete_i ;
  logic [5:0] \u_issue.u_pipe0_ctrl.mem_exception_e2_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  logic \u_issue.u_pipe0_ctrl.mul_e1_o ;
  logic \u_issue.u_pipe0_ctrl.mul_e2_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.mul_result_e2_i ;
  logic [31:0] \u_issue.u_pipe0_ctrl.opcode_e1_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.opcode_e1_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.opcode_e2_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.opcode_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.opcode_wb_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.pc_e1_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.pc_e1_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.pc_e2_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.pc_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.pc_wb_q ;
  logic [4:0] \u_issue.u_pipe0_ctrl.rd_e1_o ;
  logic [4:0] \u_issue.u_pipe0_ctrl.rd_e2_o ;
  logic [4:0] \u_issue.u_pipe0_ctrl.rd_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.result_e2_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.result_e2_q ;
  logic [31:0] \u_issue.u_pipe0_ctrl.result_e2_r ;
  logic [31:0] \u_issue.u_pipe0_ctrl.result_wb_o ;
  logic [31:0] \u_issue.u_pipe0_ctrl.result_wb_q ;
  logic \u_issue.u_pipe0_ctrl.rst_i ;
  logic \u_issue.u_pipe0_ctrl.squash_e1_e2_i ;
  logic \u_issue.u_pipe0_ctrl.squash_e1_e2_o ;
  logic \u_issue.u_pipe0_ctrl.squash_e1_e2_q ;
  logic \u_issue.u_pipe0_ctrl.squash_e1_e2_w ;
  logic \u_issue.u_pipe0_ctrl.stall_o ;
  logic \u_issue.u_pipe0_ctrl.store_e1_o ;
  logic \u_issue.u_pipe0_ctrl.take_interrupt_i ;
  logic \u_issue.u_pipe0_ctrl.valid_e1_q ;
  logic \u_issue.u_pipe0_ctrl.valid_e2_q ;
  logic \u_issue.u_pipe0_ctrl.valid_e2_w ;
  logic \u_issue.u_pipe0_ctrl.valid_wb_o ;
  logic \u_issue.u_pipe0_ctrl.valid_wb_q ;
  logic \u_issue.u_pipe1_ctrl.alu_e1_w ;
  logic [31:0] \u_issue.u_pipe1_ctrl.alu_result_e1_i ;
  logic \u_issue.u_pipe1_ctrl.branch_e1_o ;
  logic \u_issue.u_pipe1_ctrl.branch_misaligned_w ;
  logic \u_issue.u_pipe1_ctrl.clk_i ;
  logic \u_issue.u_pipe1_ctrl.csr_e1_w ;
  logic [5:0] \u_issue.u_pipe1_ctrl.csr_result_exception_e1_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.csr_result_value_e1_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.csr_result_wdata_e1_i ;
  logic \u_issue.u_pipe1_ctrl.csr_result_write_e1_i ;
  logic [11:0] \u_issue.u_pipe1_ctrl.csr_waddr_wb_o ;
  logic [9:0] \u_issue.u_pipe1_ctrl.ctrl_e1_q ;
  logic [9:0] \u_issue.u_pipe1_ctrl.ctrl_e2_q ;
  logic [9:0] \u_issue.u_pipe1_ctrl.ctrl_wb_q ;
  logic \u_issue.u_pipe1_ctrl.div_complete_i ;
  logic \u_issue.u_pipe1_ctrl.div_e1_w ;
  logic [31:0] \u_issue.u_pipe1_ctrl.div_result_i ;
  logic [5:0] \u_issue.u_pipe1_ctrl.exception_e1_q ;
  logic [5:0] \u_issue.u_pipe1_ctrl.exception_e2_q ;
  logic [5:0] \u_issue.u_pipe1_ctrl.exception_e2_r ;
  logic [5:0] \u_issue.u_pipe1_ctrl.exception_wb_o ;
  logic [5:0] \u_issue.u_pipe1_ctrl.exception_wb_q ;
  logic \u_issue.u_pipe1_ctrl.issue_accept_i ;
  logic \u_issue.u_pipe1_ctrl.issue_branch_i ;
  logic \u_issue.u_pipe1_ctrl.issue_branch_taken_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.issue_branch_target_i ;
  logic [5:0] \u_issue.u_pipe1_ctrl.issue_exception_i ;
  logic \u_issue.u_pipe1_ctrl.issue_lsu_i ;
  logic \u_issue.u_pipe1_ctrl.issue_mul_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.issue_opcode_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.issue_operand_ra_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.issue_operand_rb_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.issue_pc_i ;
  logic [4:0] \u_issue.u_pipe1_ctrl.issue_rd_i ;
  logic \u_issue.u_pipe1_ctrl.issue_rd_valid_i ;
  logic \u_issue.u_pipe1_ctrl.issue_stall_i ;
  logic \u_issue.u_pipe1_ctrl.issue_valid_i ;
  logic \u_issue.u_pipe1_ctrl.load_e1_o ;
  logic \u_issue.u_pipe1_ctrl.load_e2_o ;
  logic \u_issue.u_pipe1_ctrl.mem_complete_i ;
  logic [5:0] \u_issue.u_pipe1_ctrl.mem_exception_e2_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.mem_result_e2_i ;
  logic \u_issue.u_pipe1_ctrl.mul_e1_o ;
  logic \u_issue.u_pipe1_ctrl.mul_e2_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.mul_result_e2_i ;
  logic [31:0] \u_issue.u_pipe1_ctrl.opcode_e1_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.opcode_e1_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.opcode_e2_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.opcode_wb_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.opcode_wb_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.pc_e1_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.pc_e1_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.pc_e2_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.pc_wb_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.pc_wb_q ;
  logic [4:0] \u_issue.u_pipe1_ctrl.rd_e1_o ;
  logic [4:0] \u_issue.u_pipe1_ctrl.rd_e2_o ;
  logic [4:0] \u_issue.u_pipe1_ctrl.rd_wb_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.result_e2_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.result_e2_q ;
  logic [31:0] \u_issue.u_pipe1_ctrl.result_e2_r ;
  logic [31:0] \u_issue.u_pipe1_ctrl.result_wb_o ;
  logic [31:0] \u_issue.u_pipe1_ctrl.result_wb_q ;
  logic \u_issue.u_pipe1_ctrl.rst_i ;
  logic \u_issue.u_pipe1_ctrl.squash_e1_e2_i ;
  logic \u_issue.u_pipe1_ctrl.squash_e1_e2_o ;
  logic \u_issue.u_pipe1_ctrl.squash_e1_e2_q ;
  logic \u_issue.u_pipe1_ctrl.squash_e1_e2_w ;
  logic \u_issue.u_pipe1_ctrl.squash_wb_i ;
  logic \u_issue.u_pipe1_ctrl.stall_o ;
  logic \u_issue.u_pipe1_ctrl.store_e1_o ;
  logic \u_issue.u_pipe1_ctrl.take_interrupt_i ;
  logic \u_issue.u_pipe1_ctrl.valid_e1_q ;
  logic \u_issue.u_pipe1_ctrl.valid_e2_q ;
  logic \u_issue.u_pipe1_ctrl.valid_e2_w ;
  logic \u_issue.u_pipe1_ctrl.valid_wb_o ;
  logic \u_issue.u_pipe1_ctrl.valid_wb_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.ra0_value_r ;
  logic [31:0] \u_issue.u_regfile.REGFILE.ra1_value_r ;
  logic [31:0] \u_issue.u_regfile.REGFILE.rb0_value_r ;
  logic [31:0] \u_issue.u_regfile.REGFILE.rb1_value_r ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r10_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r11_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r12_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r13_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r14_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r15_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r16_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r17_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r18_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r19_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r1_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r20_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r21_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r22_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r23_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r24_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r25_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r26_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r27_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r28_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r29_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r2_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r30_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r31_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r3_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r4_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r5_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r6_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r7_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r8_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.reg_r9_q ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x10_a0_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x11_a1_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x12_a2_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x13_a3_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x14_a4_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x15_a5_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x16_a6_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x17_a7_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x18_s2_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x19_s3_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x1_ra_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x20_s4_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x21_s5_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x22_s6_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x23_s7_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x24_s8_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x25_s9_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x26_s10_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x27_s11_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x28_t3_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x29_t4_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x2_sp_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x30_t5_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x31_t6_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x3_gp_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x4_tp_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x5_t0_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x6_t1_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x7_t2_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x8_s0_w ;
  logic [31:0] \u_issue.u_regfile.REGFILE.x9_s1_w ;
  logic \u_issue.u_regfile.clk_i ;
  logic [4:0] \u_issue.u_regfile.ra0_i ;
  logic [31:0] \u_issue.u_regfile.ra0_value_o ;
  logic [4:0] \u_issue.u_regfile.ra1_i ;
  logic [31:0] \u_issue.u_regfile.ra1_value_o ;
  logic [4:0] \u_issue.u_regfile.rb0_i ;
  logic [31:0] \u_issue.u_regfile.rb0_value_o ;
  logic [4:0] \u_issue.u_regfile.rb1_i ;
  logic [31:0] \u_issue.u_regfile.rb1_value_o ;
  logic [4:0] \u_issue.u_regfile.rd0_i ;
  logic [31:0] \u_issue.u_regfile.rd0_value_i ;
  logic [4:0] \u_issue.u_regfile.rd1_i ;
  logic [31:0] \u_issue.u_regfile.rd1_value_i ;
  logic \u_issue.u_regfile.rst_i ;
  logic \u_issue.writeback_div_valid_i ;
  logic [31:0] \u_issue.writeback_div_value_i ;
  logic [31:0] \u_issue.writeback_exec0_value_i ;
  logic [31:0] \u_issue.writeback_exec1_value_i ;
  logic [5:0] \u_issue.writeback_mem_exception_i ;
  logic \u_issue.writeback_mem_valid_i ;
  logic [31:0] \u_issue.writeback_mem_value_i ;
  logic [31:0] \u_issue.writeback_mul_value_i ;
  logic [1:0] \u_lsu.addr_lsb_r ;
  logic \u_lsu.clk_i ;
  logic \u_lsu.complete_err_e2_w ;
  logic \u_lsu.complete_ok_e2_w ;
  logic \u_lsu.dcache_flush_w ;
  logic \u_lsu.dcache_invalidate_w ;
  logic \u_lsu.dcache_writeback_w ;
  logic \u_lsu.delay_lsu_e2_w ;
  logic \u_lsu.fault_load_align_w ;
  logic \u_lsu.fault_load_bus_w ;
  logic \u_lsu.fault_load_page_w ;
  logic \u_lsu.fault_store_align_w ;
  logic \u_lsu.fault_store_bus_w ;
  logic \u_lsu.fault_store_page_w ;
  logic \u_lsu.issue_lsu_e1_w ;
  logic \u_lsu.load_byte_r ;
  logic \u_lsu.load_half_r ;
  logic \u_lsu.load_inst_w ;
  logic \u_lsu.load_signed_inst_w ;
  logic \u_lsu.load_signed_r ;
  logic \u_lsu.mem_accept_i ;
  logic \u_lsu.mem_ack_i ;
  logic [31:0] \u_lsu.mem_addr_o ;
  logic [31:0] \u_lsu.mem_addr_q ;
  logic [31:0] \u_lsu.mem_addr_r ;
  logic \u_lsu.mem_cacheable_o ;
  logic \u_lsu.mem_cacheable_q ;
  logic [31:0] \u_lsu.mem_data_r ;
  logic [31:0] \u_lsu.mem_data_rd_i ;
  logic [31:0] \u_lsu.mem_data_wr_o ;
  logic [31:0] \u_lsu.mem_data_wr_q ;
  logic \u_lsu.mem_error_i ;
  logic \u_lsu.mem_flush_o ;
  logic \u_lsu.mem_flush_q ;
  logic \u_lsu.mem_invalidate_o ;
  logic \u_lsu.mem_invalidate_q ;
  logic \u_lsu.mem_load_q ;
  logic \u_lsu.mem_ls_q ;
  logic \u_lsu.mem_rd_o ;
  logic \u_lsu.mem_rd_q ;
  logic \u_lsu.mem_rd_r ;
  logic [10:0] \u_lsu.mem_resp_tag_i ;
  logic \u_lsu.mem_unaligned_e1_q ;
  logic \u_lsu.mem_unaligned_e2_q ;
  logic \u_lsu.mem_unaligned_r ;
  logic [3:0] \u_lsu.mem_wr_o ;
  logic [3:0] \u_lsu.mem_wr_q ;
  logic [3:0] \u_lsu.mem_wr_r ;
  logic \u_lsu.mem_writeback_o ;
  logic \u_lsu.mem_writeback_q ;
  logic \u_lsu.mem_xb_q ;
  logic \u_lsu.mem_xh_q ;
  logic [31:0] \u_lsu.opcode_opcode_i ;
  logic [31:0] \u_lsu.opcode_ra_operand_i ;
  logic [31:0] \u_lsu.opcode_rb_operand_i ;
  logic \u_lsu.opcode_valid_i ;
  logic \u_lsu.pending_lsu_e2_q ;
  logic \u_lsu.req_lb_w ;
  logic \u_lsu.req_lh_w ;
  logic \u_lsu.req_sb_w ;
  logic \u_lsu.req_sh_lh_w ;
  logic \u_lsu.req_sh_w ;
  logic \u_lsu.req_sw_lw_w ;
  logic [31:0] \u_lsu.resp_addr_w ;
  logic \u_lsu.resp_byte_w ;
  logic \u_lsu.resp_half_w ;
  logic \u_lsu.resp_load_w ;
  logic \u_lsu.resp_signed_w ;
  logic \u_lsu.rst_i ;
  logic \u_lsu.stall_o ;
  logic \u_lsu.u_lsu_request.accept_o ;
  logic \u_lsu.u_lsu_request.clk_i ;
  logic [1:0] \u_lsu.u_lsu_request.count_q ;
  logic [35:0] \u_lsu.u_lsu_request.data_in_i ;
  logic [35:0] \u_lsu.u_lsu_request.data_out_o ;
  logic \u_lsu.u_lsu_request.pop_i ;
  logic \u_lsu.u_lsu_request.push_i ;
  logic [35:0] \u_lsu.u_lsu_request.ram_q[0] ;
  logic [35:0] \u_lsu.u_lsu_request.ram_q[1] ;
  logic \u_lsu.u_lsu_request.rd_ptr_q ;
  logic \u_lsu.u_lsu_request.rst_i ;
  logic \u_lsu.u_lsu_request.valid_o ;
  logic \u_lsu.u_lsu_request.wr_ptr_q ;
  logic [31:0] \u_lsu.wb_result_r ;
  logic [5:0] \u_lsu.writeback_exception_o ;
  logic \u_lsu.writeback_valid_o ;
  logic [31:0] \u_lsu.writeback_value_o ;
  logic \u_mmu.clk_i ;
  logic \u_mmu.fetch_in_accept_o ;
  logic \u_mmu.fetch_in_error_o ;
  logic \u_mmu.fetch_in_flush_i ;
  logic [63:0] \u_mmu.fetch_in_inst_o ;
  logic [31:0] \u_mmu.fetch_in_pc_i ;
  logic \u_mmu.fetch_in_rd_i ;
  logic \u_mmu.fetch_in_valid_o ;
  logic \u_mmu.fetch_out_accept_i ;
  logic \u_mmu.fetch_out_error_i ;
  logic \u_mmu.fetch_out_flush_o ;
  logic [63:0] \u_mmu.fetch_out_inst_i ;
  logic [31:0] \u_mmu.fetch_out_pc_o ;
  logic \u_mmu.fetch_out_rd_o ;
  logic \u_mmu.fetch_out_valid_i ;
  logic \u_mmu.lsu_in_accept_o ;
  logic \u_mmu.lsu_in_ack_o ;
  logic [31:0] \u_mmu.lsu_in_addr_i ;
  logic \u_mmu.lsu_in_cacheable_i ;
  logic [31:0] \u_mmu.lsu_in_data_rd_o ;
  logic [31:0] \u_mmu.lsu_in_data_wr_i ;
  logic \u_mmu.lsu_in_error_o ;
  logic \u_mmu.lsu_in_flush_i ;
  logic \u_mmu.lsu_in_invalidate_i ;
  logic \u_mmu.lsu_in_rd_i ;
  logic [10:0] \u_mmu.lsu_in_resp_tag_o ;
  logic [3:0] \u_mmu.lsu_in_wr_i ;
  logic \u_mmu.lsu_in_writeback_i ;
  logic \u_mmu.lsu_out_accept_i ;
  logic \u_mmu.lsu_out_ack_i ;
  logic [31:0] \u_mmu.lsu_out_addr_o ;
  logic \u_mmu.lsu_out_cacheable_o ;
  logic [31:0] \u_mmu.lsu_out_data_rd_i ;
  logic [31:0] \u_mmu.lsu_out_data_wr_o ;
  logic \u_mmu.lsu_out_error_i ;
  logic \u_mmu.lsu_out_flush_o ;
  logic \u_mmu.lsu_out_invalidate_o ;
  logic \u_mmu.lsu_out_rd_o ;
  logic [10:0] \u_mmu.lsu_out_resp_tag_i ;
  logic [3:0] \u_mmu.lsu_out_wr_o ;
  logic \u_mmu.lsu_out_writeback_o ;
  logic \u_mmu.mxr_i ;
  logic \u_mmu.rst_i ;
  logic [31:0] \u_mmu.satp_i ;
  logic \u_mmu.sum_i ;
  logic \u_mul.clk_i ;
  logic \u_mul.hold_i ;
  logic \u_mul.mulhi_sel_e1_q ;
  logic \u_mul.mult_inst_w ;
  logic [63:0] \u_mul.mult_result_w ;
  logic [31:0] \u_mul.opcode_opcode_i ;
  logic [31:0] \u_mul.opcode_ra_operand_i ;
  logic [31:0] \u_mul.opcode_rb_operand_i ;
  logic \u_mul.opcode_valid_i ;
  logic [32:0] \u_mul.operand_a_e1_q ;
  logic [32:0] \u_mul.operand_a_r ;
  logic [32:0] \u_mul.operand_b_e1_q ;
  logic [32:0] \u_mul.operand_b_r ;
  logic [31:0] \u_mul.result_e2_q ;
  logic [31:0] \u_mul.result_r ;
  logic \u_mul.rst_i ;
  logic [31:0] \u_mul.writeback_value_o ;
  logic writeback_div_valid_w;
  logic [31:0] writeback_div_value_w;
  logic [31:0] writeback_exec0_value_w;
  logic [31:0] writeback_exec1_value_w;
  logic [5:0] writeback_mem_exception_w;
  logic writeback_mem_valid_w;
  logic [31:0] writeback_mem_value_w;
  logic [31:0] writeback_mul_value_w;
  assign _0128_ = 1'h0 == 1'h0;
  assign _0129_ = 1'h1 == 1'h0;
  assign _0130_ = \u_frontend.u_decode.u_fifo.wr_ptr_q == 1'h0;
  assign _0131_ = 1'h0 == 1'h1;
  assign _0132_ = 1'h1 == 1'h1;
  assign _0133_ = \u_frontend.u_decode.u_fifo.wr_ptr_q == 1'h1;
  assign _0134_ = \u_frontend.u_decode.u_fifo.rd_ptr_q == 1'h0;
  assign _0135_ = \u_frontend.u_decode.u_fifo.rd_ptr_q == 1'h1;
  assign _0136_ = \u_frontend.u_npc.branch_source_i [2] == 1'h0;
  assign _0137_ = \u_frontend.u_npc.branch_source_i [3] == 1'h0;
  assign _0138_ = \u_frontend.u_npc.branch_source_i [4] == 1'h0;
  assign _0139_ = \u_frontend.u_npc.branch_source_i [2] == 1'h1;
  assign _0140_ = \u_frontend.u_npc.branch_source_i [3] == 1'h1;
  assign _0141_ = \u_frontend.u_npc.branch_source_i [4] == 1'h1;
  assign _0142_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [0] == 1'h0;
  assign _0143_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [1] == 1'h0;
  assign _0144_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [2] == 1'h0;
  assign _0145_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [0] == 1'h0;
  assign _0146_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [1] == 1'h0;
  assign _0147_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [2] == 1'h0;
  assign _0148_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [0] == 1'h1;
  assign _0149_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [0] == 1'h1;
  assign _0150_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [1] == 1'h1;
  assign _0151_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [1] == 1'h1;
  assign _0152_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r [2] == 1'h1;
  assign _0153_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [2] == 1'h1;
  assign _0154_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [0] == 1'h0;
  assign _0155_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [1] == 1'h0;
  assign _0156_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [2] == 1'h0;
  assign _0157_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [0] == 1'h1;
  assign _0158_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [1] == 1'h1;
  assign _0159_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r [2] == 1'h1;
  assign _0160_ = \u_lsu.u_lsu_request.wr_ptr_q == 1'h0;
  assign _0161_ = \u_lsu.u_lsu_request.wr_ptr_q == 1'h1;
  assign _0000_ = _0128_ & _0128_;
  assign _0001_ = _0128_ & _0000_;
  assign _0002_ = _0129_ & _0000_;
  assign _0003_ = _0129_ & _0128_;
  assign _0004_ = _0128_ & _0003_;
  assign _0005_ = _0129_ & _0003_;
  assign _0006_ = _0128_ & _0129_;
  assign _0007_ = _0128_ & _0006_;
  assign _0008_ = _0129_ & _0006_;
  assign _0009_ = _0129_ & _0129_;
  assign _0010_ = _0128_ & _0009_;
  assign _0011_ = _0129_ & _0009_;
  assign _0012_ = _0137_ & _0138_;
  assign _0013_ = _0136_ & _0012_;
  assign _0014_ = _0131_ & _0000_;
  assign _0015_ = _0132_ & _0000_;
  assign _0016_ = _0131_ & _0003_;
  assign _0017_ = _0132_ & _0003_;
  assign _0018_ = _0131_ & _0006_;
  assign _0019_ = _0132_ & _0006_;
  assign _0020_ = _0131_ & _0009_;
  assign _0021_ = _0132_ & _0009_;
  assign _0022_ = _0139_ & _0012_;
  assign _0023_ = _0131_ & _0128_;
  assign _0024_ = _0128_ & _0023_;
  assign _0025_ = _0129_ & _0023_;
  assign _0026_ = _0132_ & _0128_;
  assign _0027_ = _0128_ & _0026_;
  assign _0028_ = _0129_ & _0026_;
  assign _0029_ = _0131_ & _0129_;
  assign _0030_ = _0128_ & _0029_;
  assign _0031_ = _0129_ & _0029_;
  assign _0032_ = _0132_ & _0129_;
  assign _0033_ = _0128_ & _0032_;
  assign _0034_ = _0129_ & _0032_;
  assign _0035_ = _0140_ & _0138_;
  assign _0036_ = _0136_ & _0035_;
  assign _0037_ = _0131_ & _0023_;
  assign _0038_ = _0132_ & _0023_;
  assign _0039_ = _0131_ & _0026_;
  assign _0040_ = _0132_ & _0026_;
  assign _0041_ = _0131_ & _0029_;
  assign _0042_ = _0132_ & _0029_;
  assign _0043_ = _0131_ & _0032_;
  assign _0044_ = _0132_ & _0032_;
  assign _0045_ = _0139_ & _0035_;
  assign _0046_ = _0128_ & _0131_;
  assign _0047_ = _0128_ & _0046_;
  assign _0048_ = _0129_ & _0046_;
  assign _0049_ = _0129_ & _0131_;
  assign _0050_ = _0128_ & _0049_;
  assign _0051_ = _0129_ & _0049_;
  assign _0052_ = _0128_ & _0132_;
  assign _0053_ = _0128_ & _0052_;
  assign _0054_ = _0129_ & _0052_;
  assign _0055_ = _0129_ & _0132_;
  assign _0056_ = _0128_ & _0055_;
  assign _0057_ = _0129_ & _0055_;
  assign _0058_ = _0137_ & _0141_;
  assign _0059_ = _0136_ & _0058_;
  assign _0060_ = _0131_ & _0046_;
  assign _0061_ = _0132_ & _0046_;
  assign _0062_ = _0131_ & _0049_;
  assign _0063_ = _0132_ & _0049_;
  assign _0064_ = _0131_ & _0052_;
  assign _0065_ = _0132_ & _0052_;
  assign _0066_ = _0131_ & _0055_;
  assign _0067_ = _0132_ & _0055_;
  assign _0068_ = _0139_ & _0058_;
  assign _0069_ = _0131_ & _0131_;
  assign _0070_ = _0128_ & _0069_;
  assign _0071_ = _0129_ & _0069_;
  assign _0072_ = _0132_ & _0131_;
  assign _0073_ = _0128_ & _0072_;
  assign _0074_ = _0129_ & _0072_;
  assign _0075_ = _0131_ & _0132_;
  assign _0076_ = _0128_ & _0075_;
  assign _0077_ = _0129_ & _0075_;
  assign _0078_ = _0132_ & _0132_;
  assign _0079_ = _0128_ & _0078_;
  assign _0080_ = _0129_ & _0078_;
  assign _0081_ = _0140_ & _0141_;
  assign _0082_ = _0136_ & _0081_;
  assign _0083_ = _0131_ & _0069_;
  assign _0084_ = _0132_ & _0069_;
  assign _0085_ = _0131_ & _0072_;
  assign _0086_ = _0132_ & _0072_;
  assign _0087_ = _0131_ & _0075_;
  assign _0088_ = _0132_ & _0075_;
  assign _0089_ = _0131_ & _0078_;
  assign _0090_ = _0132_ & _0078_;
  assign _0091_ = _0139_ & _0081_;
  assign _0092_ = _0143_ & _0144_;
  assign _0093_ = _0142_ & _0092_;
  assign _0094_ = _0146_ & _0147_;
  assign _0095_ = _0145_ & _0094_;
  assign _0096_ = _0148_ & _0092_;
  assign _0097_ = _0149_ & _0094_;
  assign _0098_ = _0150_ & _0144_;
  assign _0099_ = _0142_ & _0098_;
  assign _0100_ = _0151_ & _0147_;
  assign _0101_ = _0145_ & _0100_;
  assign _0102_ = _0148_ & _0098_;
  assign _0103_ = _0149_ & _0100_;
  assign _0104_ = _0143_ & _0152_;
  assign _0105_ = _0142_ & _0104_;
  assign _0106_ = _0146_ & _0153_;
  assign _0107_ = _0145_ & _0106_;
  assign _0108_ = _0148_ & _0104_;
  assign _0109_ = _0149_ & _0106_;
  assign _0110_ = _0150_ & _0152_;
  assign _0111_ = _0142_ & _0110_;
  assign _0112_ = _0151_ & _0153_;
  assign _0113_ = _0145_ & _0112_;
  assign _0114_ = _0148_ & _0110_;
  assign _0115_ = _0149_ & _0112_;
  assign _0116_ = _0155_ & _0156_;
  assign _0117_ = _0154_ & _0116_;
  assign _0118_ = _0157_ & _0116_;
  assign _0119_ = _0158_ & _0156_;
  assign _0120_ = _0154_ & _0119_;
  assign _0121_ = _0157_ & _0119_;
  assign _0122_ = _0155_ & _0159_;
  assign _0123_ = _0154_ & _0122_;
  assign _0124_ = _0157_ & _0122_;
  assign _0125_ = _0158_ & _0159_;
  assign _0126_ = _0154_ & _0125_;
  assign _0127_ = _0157_ & _0125_;
  assign \u_frontend.u_decode.u_fifo.info0_out_o = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.info0_q[1] : \u_frontend.u_decode.u_fifo.info0_q[0] ;
  assign _0162_ = _0128_ & _2739_[1];
  assign _0163_ = _0129_ & _2739_[1];
  assign _0164_ = _0128_ & _2740_[1];
  assign _0165_ = _0129_ & _2740_[1];
  assign _0166_ = _0130_ & _2741_[1];
  assign _0167_ = _0131_ & _2739_[1];
  assign _0168_ = _0132_ & _2739_[1];
  assign _0169_ = _0131_ & _2740_[1];
  assign _0170_ = _0132_ & _2740_[1];
  assign _0171_ = _0133_ & _2741_[1];
  assign _0172_ = _0162_ ? 2'h0 : \u_frontend.u_decode.u_fifo.info0_q[0] ;
  assign _0173_ = _0163_ ? 2'h0 : _0172_;
  assign _0174_ = _0164_ ? 2'h0 : _0173_;
  assign _0175_ = _0165_ ? 2'h0 : _0174_;
  logic [1:0] fangyuan0;
  assign fangyuan0 = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign _0176_ = _0166_ ? fangyuan0 : _0175_;
  assign _0177_ = _0167_ ? 2'h0 : \u_frontend.u_decode.u_fifo.info0_q[1] ;
  assign _0178_ = _0168_ ? 2'h0 : _0177_;
  assign _0179_ = _0169_ ? 2'h0 : _0178_;
  assign _0180_ = _0170_ ? 2'h0 : _0179_;
  logic [1:0] fangyuan1;
  assign fangyuan1 = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign _0181_ = _0171_ ? fangyuan1 : _0180_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.info0_q[0] <= _0176_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.info0_q[1] <= _0181_;
  assign \u_frontend.u_decode.u_fifo.info1_out_o = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.info1_q[1] : \u_frontend.u_decode.u_fifo.info1_q[0] ;
  assign _0182_ = _0128_ & _2739_[1];
  assign _0183_ = _0129_ & _2739_[1];
  assign _0184_ = _0128_ & _2740_[1];
  assign _0185_ = _0129_ & _2740_[1];
  assign _0186_ = _0130_ & _2741_[1];
  assign _0187_ = _0131_ & _2739_[1];
  assign _0188_ = _0132_ & _2739_[1];
  assign _0189_ = _0131_ & _2740_[1];
  assign _0190_ = _0132_ & _2740_[1];
  assign _0191_ = _0133_ & _2741_[1];
  assign _0192_ = _0182_ ? 2'h0 : \u_frontend.u_decode.u_fifo.info1_q[0] ;
  assign _0193_ = _0183_ ? 2'h0 : _0192_;
  assign _0194_ = _0184_ ? 2'h0 : _0193_;
  assign _0195_ = _0185_ ? 2'h0 : _0194_;
  logic [1:0] fangyuan2;
  assign fangyuan2 = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign _0196_ = _0186_ ? fangyuan2 : _0195_;
  assign _0197_ = _0187_ ? 2'h0 : \u_frontend.u_decode.u_fifo.info1_q[1] ;
  assign _0198_ = _0188_ ? 2'h0 : _0197_;
  assign _0199_ = _0189_ ? 2'h0 : _0198_;
  assign _0200_ = _0190_ ? 2'h0 : _0199_;
  logic [1:0] fangyuan3;
  assign fangyuan3 = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign _0201_ = _0191_ ? fangyuan3 : _0200_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.info1_q[0] <= _0196_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.info1_q[1] <= _0201_;
  logic [31:0] fangyuan4;
  assign { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], _2738_ } = fangyuan4;
  assign fangyuan4 = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.pc_q[1] : \u_frontend.u_decode.u_fifo.pc_q[0] ;
  assign _0202_ = _0128_ & _2739_[1];
  assign _0203_ = _0129_ & _2739_[1];
  assign _0204_ = _0130_ & _2741_[1];
  assign _0205_ = _0131_ & _2739_[1];
  assign _0206_ = _0132_ & _2739_[1];
  assign _0207_ = _0133_ & _2741_[1];
  assign _0208_ = _0202_ ? 32'h00000000 : \u_frontend.u_decode.u_fifo.pc_q[0] ;
  assign _0209_ = _0203_ ? 32'h00000000 : _0208_;
  assign _0210_ = _0204_ ? \u_frontend.u_decode.u_fifo.pc_in_i : _0209_;
  assign _0211_ = _0205_ ? 32'h00000000 : \u_frontend.u_decode.u_fifo.pc_q[1] ;
  assign _0212_ = _0206_ ? 32'h00000000 : _0211_;
  assign _0213_ = _0207_ ? \u_frontend.u_decode.u_fifo.pc_in_i : _0212_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.pc_q[0] <= _0210_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.pc_q[1] <= _0213_;
  logic [63:0] fangyuan5;
  assign { \u_frontend.u_decode.u_fifo.data1_out_o , \u_frontend.u_decode.u_fifo.data0_out_o } = fangyuan5;
  assign fangyuan5 = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.ram_q[1] : \u_frontend.u_decode.u_fifo.ram_q[0] ;
  assign _0214_ = _0128_ & _2739_[1];
  assign _0215_ = _0129_ & _2739_[1];
  assign _0216_ = _0130_ & _2741_[1];
  assign _0217_ = _0131_ & _2739_[1];
  assign _0218_ = _0132_ & _2739_[1];
  assign _0219_ = _0133_ & _2741_[1];
  assign _0220_ = _0214_ ? 64'h0000000000000000 : \u_frontend.u_decode.u_fifo.ram_q[0] ;
  assign _0221_ = _0215_ ? 64'h0000000000000000 : _0220_;
  assign _0222_ = _0216_ ? \u_frontend.u_decode.u_fifo.data_in_i : _0221_;
  assign _0223_ = _0217_ ? 64'h0000000000000000 : \u_frontend.u_decode.u_fifo.ram_q[1] ;
  assign _0224_ = _0218_ ? 64'h0000000000000000 : _0223_;
  assign _0225_ = _0219_ ? \u_frontend.u_decode.u_fifo.data_in_i : _0224_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.ram_q[0] <= _0222_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.ram_q[1] <= _0225_;
  assign _2757_ = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.valid0_q[1] : \u_frontend.u_decode.u_fifo.valid0_q[0] ;
  assign _0226_ = _0128_ & _2739_[1];
  assign _0227_ = _0129_ & _2739_[1];
  assign _0228_ = _0130_ & _2741_[1];
  assign _0229_ = _0134_ & _2742_;
  assign _0230_ = _0131_ & _2739_[1];
  assign _0231_ = _0132_ & _2739_[1];
  assign _0232_ = _0133_ & _2741_[1];
  assign _0233_ = _0135_ & _2742_;
  assign _0234_ = _0226_ ? 1'h0 : \u_frontend.u_decode.u_fifo.valid0_q[0] ;
  assign _0235_ = _0227_ ? 1'h0 : _0234_;
  assign _0236_ = _0228_ ? 1'h1 : _0235_;
  assign _0237_ = _0229_ ? 1'h0 : _0236_;
  assign _0238_ = _0230_ ? 1'h0 : \u_frontend.u_decode.u_fifo.valid0_q[1] ;
  assign _0239_ = _0231_ ? 1'h0 : _0238_;
  assign _0240_ = _0232_ ? 1'h1 : _0239_;
  assign _0241_ = _0233_ ? 1'h0 : _0240_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.valid0_q[0] <= _0237_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.valid0_q[1] <= _0241_;
  assign _2758_ = \u_frontend.u_decode.u_fifo.rd_ptr_q ? \u_frontend.u_decode.u_fifo.valid1_q[1] : \u_frontend.u_decode.u_fifo.valid1_q[0] ;
  assign _0242_ = _0128_ & _2739_[1];
  assign _0243_ = _0129_ & _2739_[1];
  assign _0244_ = _0130_ & _2741_[1];
  assign _0245_ = _0134_ & _2744_;
  assign _0246_ = _0131_ & _2739_[1];
  assign _0247_ = _0132_ & _2739_[1];
  assign _0248_ = _0133_ & _2741_[1];
  assign _0249_ = _0135_ & _2744_;
  assign _0250_ = _0242_ ? 1'h0 : \u_frontend.u_decode.u_fifo.valid1_q[0] ;
  assign _0251_ = _0243_ ? 1'h0 : _0250_;
  assign _0252_ = _0244_ ? _2743_ : _0251_;
  assign _0253_ = _0245_ ? 1'h0 : _0252_;
  assign _0254_ = _0246_ ? 1'h0 : \u_frontend.u_decode.u_fifo.valid1_q[1] ;
  assign _0255_ = _0247_ ? 1'h0 : _0254_;
  assign _0256_ = _0248_ ? _2743_ : _0255_;
  assign _0257_ = _0249_ ? 1'h0 : _0256_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.valid1_q[0] <= _0253_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.valid1_q[1] <= _0257_;
  assign _2999_ = \u_frontend.u_npc.branch_source_i [4] ? _0259_ : _0258_;
  assign _0258_ = \u_frontend.u_npc.branch_source_i [3] ? _0261_ : _0260_;
  assign _0259_ = \u_frontend.u_npc.branch_source_i [3] ? _0263_ : _0262_;
  assign _0260_ = \u_frontend.u_npc.branch_source_i [2] ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[0] ;
  assign _0261_ = \u_frontend.u_npc.branch_source_i [2] ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[2] ;
  assign _0262_ = \u_frontend.u_npc.branch_source_i [2] ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[4] ;
  assign _0263_ = \u_frontend.u_npc.branch_source_i [2] ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[6] ;
  assign _3000_ = \u_frontend.u_fetch.icache_pc_w [4] ? _0265_ : _0264_;
  assign _0264_ = \u_frontend.u_fetch.icache_pc_w [3] ? _0267_ : _0266_;
  assign _0265_ = \u_frontend.u_fetch.icache_pc_w [3] ? _0269_ : _0268_;
  assign _0266_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[0] ;
  assign _0267_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[2] ;
  assign _0268_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[4] ;
  assign _0269_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ? \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[6] ;
  assign _0270_ = _0001_ & _2827_[1];
  assign _0271_ = _0002_ & _2827_[1];
  assign _0272_ = _0004_ & _2827_[1];
  assign _0273_ = _0005_ & _2827_[1];
  assign _0274_ = _0007_ & _2827_[1];
  assign _0275_ = _0008_ & _2827_[1];
  assign _0276_ = _0010_ & _2827_[1];
  assign _0277_ = _0011_ & _2827_[1];
  assign _0278_ = _0013_ & _2829_[1];
  assign _0279_ = _0013_ & _2831_[1];
  assign _0280_ = _0014_ & _2827_[1];
  assign _0281_ = _0015_ & _2827_[1];
  assign _0282_ = _0016_ & _2827_[1];
  assign _0283_ = _0017_ & _2827_[1];
  assign _0284_ = _0018_ & _2827_[1];
  assign _0285_ = _0019_ & _2827_[1];
  assign _0286_ = _0020_ & _2827_[1];
  assign _0287_ = _0021_ & _2827_[1];
  assign _0288_ = _0022_ & _2829_[1];
  assign _0289_ = _0022_ & _2831_[1];
  assign _0290_ = _0024_ & _2827_[1];
  assign _0291_ = _0025_ & _2827_[1];
  assign _0292_ = _0027_ & _2827_[1];
  assign _0293_ = _0028_ & _2827_[1];
  assign _0294_ = _0030_ & _2827_[1];
  assign _0295_ = _0031_ & _2827_[1];
  assign _0296_ = _0033_ & _2827_[1];
  assign _0297_ = _0034_ & _2827_[1];
  assign _0298_ = _0036_ & _2829_[1];
  assign _0299_ = _0036_ & _2831_[1];
  assign _0300_ = _0037_ & _2827_[1];
  assign _0301_ = _0038_ & _2827_[1];
  assign _0302_ = _0039_ & _2827_[1];
  assign _0303_ = _0040_ & _2827_[1];
  assign _0304_ = _0041_ & _2827_[1];
  assign _0305_ = _0042_ & _2827_[1];
  assign _0306_ = _0043_ & _2827_[1];
  assign _0307_ = _0044_ & _2827_[1];
  assign _0308_ = _0045_ & _2829_[1];
  assign _0309_ = _0045_ & _2831_[1];
  assign _0310_ = _0047_ & _2827_[1];
  assign _0311_ = _0048_ & _2827_[1];
  assign _0312_ = _0050_ & _2827_[1];
  assign _0313_ = _0051_ & _2827_[1];
  assign _0314_ = _0053_ & _2827_[1];
  assign _0315_ = _0054_ & _2827_[1];
  assign _0316_ = _0056_ & _2827_[1];
  assign _0317_ = _0057_ & _2827_[1];
  assign _0318_ = _0059_ & _2829_[1];
  assign _0319_ = _0059_ & _2831_[1];
  assign _0320_ = _0060_ & _2827_[1];
  assign _0321_ = _0061_ & _2827_[1];
  assign _0322_ = _0062_ & _2827_[1];
  assign _0323_ = _0063_ & _2827_[1];
  assign _0324_ = _0064_ & _2827_[1];
  assign _0325_ = _0065_ & _2827_[1];
  assign _0326_ = _0066_ & _2827_[1];
  assign _0327_ = _0067_ & _2827_[1];
  assign _0328_ = _0068_ & _2829_[1];
  assign _0329_ = _0068_ & _2831_[1];
  assign _0330_ = _0070_ & _2827_[1];
  assign _0331_ = _0071_ & _2827_[1];
  assign _0332_ = _0073_ & _2827_[1];
  assign _0333_ = _0074_ & _2827_[1];
  assign _0334_ = _0076_ & _2827_[1];
  assign _0335_ = _0077_ & _2827_[1];
  assign _0336_ = _0079_ & _2827_[1];
  assign _0337_ = _0080_ & _2827_[1];
  assign _0338_ = _0082_ & _2829_[1];
  assign _0339_ = _0082_ & _2831_[1];
  assign _0340_ = _0083_ & _2827_[1];
  assign _0341_ = _0084_ & _2827_[1];
  assign _0342_ = _0085_ & _2827_[1];
  assign _0343_ = _0086_ & _2827_[1];
  assign _0344_ = _0087_ & _2827_[1];
  assign _0345_ = _0088_ & _2827_[1];
  assign _0346_ = _0089_ & _2827_[1];
  assign _0347_ = _0090_ & _2827_[1];
  assign _0348_ = _0091_ & _2829_[1];
  assign _0349_ = _0091_ & _2831_[1];
  assign _0350_ = _0270_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[0] ;
  assign _0351_ = _0271_ ? 2'h3 : _0350_;
  assign _0352_ = _0272_ ? 2'h3 : _0351_;
  assign _0353_ = _0273_ ? 2'h3 : _0352_;
  assign _0354_ = _0274_ ? 2'h3 : _0353_;
  assign _0355_ = _0275_ ? 2'h3 : _0354_;
  assign _0356_ = _0276_ ? 2'h3 : _0355_;
  assign _0357_ = _0277_ ? 2'h3 : _0356_;
  assign _0358_ = _0278_ ? _2828_ : _0357_;
  assign _0359_ = _0279_ ? _2830_ : _0358_;
  assign _0360_ = _0280_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[1] ;
  assign _0361_ = _0281_ ? 2'h3 : _0360_;
  assign _0362_ = _0282_ ? 2'h3 : _0361_;
  assign _0363_ = _0283_ ? 2'h3 : _0362_;
  assign _0364_ = _0284_ ? 2'h3 : _0363_;
  assign _0365_ = _0285_ ? 2'h3 : _0364_;
  assign _0366_ = _0286_ ? 2'h3 : _0365_;
  assign _0367_ = _0287_ ? 2'h3 : _0366_;
  assign _0368_ = _0288_ ? _2828_ : _0367_;
  assign _0369_ = _0289_ ? _2830_ : _0368_;
  assign _0370_ = _0290_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[2] ;
  assign _0371_ = _0291_ ? 2'h3 : _0370_;
  assign _0372_ = _0292_ ? 2'h3 : _0371_;
  assign _0373_ = _0293_ ? 2'h3 : _0372_;
  assign _0374_ = _0294_ ? 2'h3 : _0373_;
  assign _0375_ = _0295_ ? 2'h3 : _0374_;
  assign _0376_ = _0296_ ? 2'h3 : _0375_;
  assign _0377_ = _0297_ ? 2'h3 : _0376_;
  assign _0378_ = _0298_ ? _2828_ : _0377_;
  assign _0379_ = _0299_ ? _2830_ : _0378_;
  assign _0380_ = _0300_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[3] ;
  assign _0381_ = _0301_ ? 2'h3 : _0380_;
  assign _0382_ = _0302_ ? 2'h3 : _0381_;
  assign _0383_ = _0303_ ? 2'h3 : _0382_;
  assign _0384_ = _0304_ ? 2'h3 : _0383_;
  assign _0385_ = _0305_ ? 2'h3 : _0384_;
  assign _0386_ = _0306_ ? 2'h3 : _0385_;
  assign _0387_ = _0307_ ? 2'h3 : _0386_;
  assign _0388_ = _0308_ ? _2828_ : _0387_;
  assign _0389_ = _0309_ ? _2830_ : _0388_;
  assign _0390_ = _0310_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[4] ;
  assign _0391_ = _0311_ ? 2'h3 : _0390_;
  assign _0392_ = _0312_ ? 2'h3 : _0391_;
  assign _0393_ = _0313_ ? 2'h3 : _0392_;
  assign _0394_ = _0314_ ? 2'h3 : _0393_;
  assign _0395_ = _0315_ ? 2'h3 : _0394_;
  assign _0396_ = _0316_ ? 2'h3 : _0395_;
  assign _0397_ = _0317_ ? 2'h3 : _0396_;
  assign _0398_ = _0318_ ? _2828_ : _0397_;
  assign _0399_ = _0319_ ? _2830_ : _0398_;
  assign _0400_ = _0320_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[5] ;
  assign _0401_ = _0321_ ? 2'h3 : _0400_;
  assign _0402_ = _0322_ ? 2'h3 : _0401_;
  assign _0403_ = _0323_ ? 2'h3 : _0402_;
  assign _0404_ = _0324_ ? 2'h3 : _0403_;
  assign _0405_ = _0325_ ? 2'h3 : _0404_;
  assign _0406_ = _0326_ ? 2'h3 : _0405_;
  assign _0407_ = _0327_ ? 2'h3 : _0406_;
  assign _0408_ = _0328_ ? _2828_ : _0407_;
  assign _0409_ = _0329_ ? _2830_ : _0408_;
  assign _0410_ = _0330_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[6] ;
  assign _0411_ = _0331_ ? 2'h3 : _0410_;
  assign _0412_ = _0332_ ? 2'h3 : _0411_;
  assign _0413_ = _0333_ ? 2'h3 : _0412_;
  assign _0414_ = _0334_ ? 2'h3 : _0413_;
  assign _0415_ = _0335_ ? 2'h3 : _0414_;
  assign _0416_ = _0336_ ? 2'h3 : _0415_;
  assign _0417_ = _0337_ ? 2'h3 : _0416_;
  assign _0418_ = _0338_ ? _2828_ : _0417_;
  assign _0419_ = _0339_ ? _2830_ : _0418_;
  assign _0420_ = _0340_ ? 2'h3 : \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[7] ;
  assign _0421_ = _0341_ ? 2'h3 : _0420_;
  assign _0422_ = _0342_ ? 2'h3 : _0421_;
  assign _0423_ = _0343_ ? 2'h3 : _0422_;
  assign _0424_ = _0344_ ? 2'h3 : _0423_;
  assign _0425_ = _0345_ ? 2'h3 : _0424_;
  assign _0426_ = _0346_ ? 2'h3 : _0425_;
  assign _0427_ = _0347_ ? 2'h3 : _0426_;
  assign _0428_ = _0348_ ? _2828_ : _0427_;
  assign _0429_ = _0349_ ? _2830_ : _0428_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[0] <= _0359_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[1] <= _0369_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[2] <= _0379_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[3] <= _0389_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[4] <= _0399_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[5] <= _0409_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[6] <= _0419_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.bht_sat_q[7] <= _0429_;
  assign _3001_ = 1'h0 ? _0431_ : _0430_;
  assign _0430_ = 1'h0 ? _0433_ : _0432_;
  assign _0431_ = 1'h0 ? _0435_ : _0434_;
  assign _0432_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0433_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0434_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0435_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3002_ = 1'h0 ? _0437_ : _0436_;
  assign _0436_ = 1'h0 ? _0439_ : _0438_;
  assign _0437_ = 1'h0 ? _0441_ : _0440_;
  assign _0438_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0439_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0440_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0441_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3003_ = 1'h0 ? _0443_ : _0442_;
  assign _0442_ = 1'h1 ? _0445_ : _0444_;
  assign _0443_ = 1'h1 ? _0447_ : _0446_;
  assign _0444_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0445_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0446_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0447_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3004_ = 1'h0 ? _0449_ : _0448_;
  assign _0448_ = 1'h1 ? _0451_ : _0450_;
  assign _0449_ = 1'h1 ? _0453_ : _0452_;
  assign _0450_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0451_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0452_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0453_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3005_ = 1'h1 ? _0455_ : _0454_;
  assign _0454_ = 1'h0 ? _0457_ : _0456_;
  assign _0455_ = 1'h0 ? _0459_ : _0458_;
  assign _0456_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0457_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0458_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0459_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3006_ = 1'h1 ? _0461_ : _0460_;
  assign _0460_ = 1'h0 ? _0463_ : _0462_;
  assign _0461_ = 1'h0 ? _0465_ : _0464_;
  assign _0462_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0463_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0464_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0465_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3007_ = 1'h1 ? _0467_ : _0466_;
  assign _0466_ = 1'h1 ? _0469_ : _0468_;
  assign _0467_ = 1'h1 ? _0471_ : _0470_;
  assign _0468_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0469_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0470_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0471_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _3008_ = 1'h1 ? _0473_ : _0472_;
  assign _0472_ = 1'h1 ? _0475_ : _0474_;
  assign _0473_ = 1'h1 ? _0477_ : _0476_;
  assign _0474_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0475_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0476_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0477_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _0478_ = _0001_ & _2827_[1];
  assign _0479_ = _0002_ & _2827_[1];
  assign _0480_ = _0004_ & _2827_[1];
  assign _0481_ = _0005_ & _2827_[1];
  assign _0482_ = _0007_ & _2827_[1];
  assign _0483_ = _0008_ & _2827_[1];
  assign _0484_ = _0010_ & _2827_[1];
  assign _0485_ = _0011_ & _2827_[1];
  assign _0486_ = _0093_ & _2832_;
  assign _0487_ = _0095_ & _2833_;
  assign _0488_ = _0014_ & _2827_[1];
  assign _0489_ = _0015_ & _2827_[1];
  assign _0490_ = _0016_ & _2827_[1];
  assign _0491_ = _0017_ & _2827_[1];
  assign _0492_ = _0018_ & _2827_[1];
  assign _0493_ = _0019_ & _2827_[1];
  assign _0494_ = _0020_ & _2827_[1];
  assign _0495_ = _0021_ & _2827_[1];
  assign _0496_ = _0096_ & _2832_;
  assign _0497_ = _0097_ & _2833_;
  assign _0498_ = _0024_ & _2827_[1];
  assign _0499_ = _0025_ & _2827_[1];
  assign _0500_ = _0027_ & _2827_[1];
  assign _0501_ = _0028_ & _2827_[1];
  assign _0502_ = _0030_ & _2827_[1];
  assign _0503_ = _0031_ & _2827_[1];
  assign _0504_ = _0033_ & _2827_[1];
  assign _0505_ = _0034_ & _2827_[1];
  assign _0506_ = _0099_ & _2832_;
  assign _0507_ = _0101_ & _2833_;
  assign _0508_ = _0037_ & _2827_[1];
  assign _0509_ = _0038_ & _2827_[1];
  assign _0510_ = _0039_ & _2827_[1];
  assign _0511_ = _0040_ & _2827_[1];
  assign _0512_ = _0041_ & _2827_[1];
  assign _0513_ = _0042_ & _2827_[1];
  assign _0514_ = _0043_ & _2827_[1];
  assign _0515_ = _0044_ & _2827_[1];
  assign _0516_ = _0102_ & _2832_;
  assign _0517_ = _0103_ & _2833_;
  assign _0518_ = _0047_ & _2827_[1];
  assign _0519_ = _0048_ & _2827_[1];
  assign _0520_ = _0050_ & _2827_[1];
  assign _0521_ = _0051_ & _2827_[1];
  assign _0522_ = _0053_ & _2827_[1];
  assign _0523_ = _0054_ & _2827_[1];
  assign _0524_ = _0056_ & _2827_[1];
  assign _0525_ = _0057_ & _2827_[1];
  assign _0526_ = _0105_ & _2832_;
  assign _0527_ = _0107_ & _2833_;
  assign _0528_ = _0060_ & _2827_[1];
  assign _0529_ = _0061_ & _2827_[1];
  assign _0530_ = _0062_ & _2827_[1];
  assign _0531_ = _0063_ & _2827_[1];
  assign _0532_ = _0064_ & _2827_[1];
  assign _0533_ = _0065_ & _2827_[1];
  assign _0534_ = _0066_ & _2827_[1];
  assign _0535_ = _0067_ & _2827_[1];
  assign _0536_ = _0108_ & _2832_;
  assign _0537_ = _0109_ & _2833_;
  assign _0538_ = _0070_ & _2827_[1];
  assign _0539_ = _0071_ & _2827_[1];
  assign _0540_ = _0073_ & _2827_[1];
  assign _0541_ = _0074_ & _2827_[1];
  assign _0542_ = _0076_ & _2827_[1];
  assign _0543_ = _0077_ & _2827_[1];
  assign _0544_ = _0079_ & _2827_[1];
  assign _0545_ = _0080_ & _2827_[1];
  assign _0546_ = _0111_ & _2832_;
  assign _0547_ = _0113_ & _2833_;
  assign _0548_ = _0083_ & _2827_[1];
  assign _0549_ = _0084_ & _2827_[1];
  assign _0550_ = _0085_ & _2827_[1];
  assign _0551_ = _0086_ & _2827_[1];
  assign _0552_ = _0087_ & _2827_[1];
  assign _0553_ = _0088_ & _2827_[1];
  assign _0554_ = _0089_ & _2827_[1];
  assign _0555_ = _0090_ & _2827_[1];
  assign _0556_ = _0114_ & _2832_;
  assign _0557_ = _0115_ & _2833_;
  assign _0558_ = _0478_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] ;
  assign _0559_ = _0479_ ? 1'h0 : _0558_;
  assign _0560_ = _0480_ ? 1'h0 : _0559_;
  assign _0561_ = _0481_ ? 1'h0 : _0560_;
  assign _0562_ = _0482_ ? 1'h0 : _0561_;
  assign _0563_ = _0483_ ? 1'h0 : _0562_;
  assign _0564_ = _0484_ ? 1'h0 : _0563_;
  assign _0565_ = _0485_ ? 1'h0 : _0564_;
  assign _0566_ = _0486_ ? \u_frontend.u_npc.branch_is_call_i : _0565_;
  assign _0567_ = _0487_ ? \u_frontend.u_npc.branch_is_call_i : _0566_;
  assign _0568_ = _0488_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] ;
  assign _0569_ = _0489_ ? 1'h0 : _0568_;
  assign _0570_ = _0490_ ? 1'h0 : _0569_;
  assign _0571_ = _0491_ ? 1'h0 : _0570_;
  assign _0572_ = _0492_ ? 1'h0 : _0571_;
  assign _0573_ = _0493_ ? 1'h0 : _0572_;
  assign _0574_ = _0494_ ? 1'h0 : _0573_;
  assign _0575_ = _0495_ ? 1'h0 : _0574_;
  assign _0576_ = _0496_ ? \u_frontend.u_npc.branch_is_call_i : _0575_;
  assign _0577_ = _0497_ ? \u_frontend.u_npc.branch_is_call_i : _0576_;
  assign _0578_ = _0498_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] ;
  assign _0579_ = _0499_ ? 1'h0 : _0578_;
  assign _0580_ = _0500_ ? 1'h0 : _0579_;
  assign _0581_ = _0501_ ? 1'h0 : _0580_;
  assign _0582_ = _0502_ ? 1'h0 : _0581_;
  assign _0583_ = _0503_ ? 1'h0 : _0582_;
  assign _0584_ = _0504_ ? 1'h0 : _0583_;
  assign _0585_ = _0505_ ? 1'h0 : _0584_;
  assign _0586_ = _0506_ ? \u_frontend.u_npc.branch_is_call_i : _0585_;
  assign _0587_ = _0507_ ? \u_frontend.u_npc.branch_is_call_i : _0586_;
  assign _0588_ = _0508_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] ;
  assign _0589_ = _0509_ ? 1'h0 : _0588_;
  assign _0590_ = _0510_ ? 1'h0 : _0589_;
  assign _0591_ = _0511_ ? 1'h0 : _0590_;
  assign _0592_ = _0512_ ? 1'h0 : _0591_;
  assign _0593_ = _0513_ ? 1'h0 : _0592_;
  assign _0594_ = _0514_ ? 1'h0 : _0593_;
  assign _0595_ = _0515_ ? 1'h0 : _0594_;
  assign _0596_ = _0516_ ? \u_frontend.u_npc.branch_is_call_i : _0595_;
  assign _0597_ = _0517_ ? \u_frontend.u_npc.branch_is_call_i : _0596_;
  assign _0598_ = _0518_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] ;
  assign _0599_ = _0519_ ? 1'h0 : _0598_;
  assign _0600_ = _0520_ ? 1'h0 : _0599_;
  assign _0601_ = _0521_ ? 1'h0 : _0600_;
  assign _0602_ = _0522_ ? 1'h0 : _0601_;
  assign _0603_ = _0523_ ? 1'h0 : _0602_;
  assign _0604_ = _0524_ ? 1'h0 : _0603_;
  assign _0605_ = _0525_ ? 1'h0 : _0604_;
  assign _0606_ = _0526_ ? \u_frontend.u_npc.branch_is_call_i : _0605_;
  assign _0607_ = _0527_ ? \u_frontend.u_npc.branch_is_call_i : _0606_;
  assign _0608_ = _0528_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] ;
  assign _0609_ = _0529_ ? 1'h0 : _0608_;
  assign _0610_ = _0530_ ? 1'h0 : _0609_;
  assign _0611_ = _0531_ ? 1'h0 : _0610_;
  assign _0612_ = _0532_ ? 1'h0 : _0611_;
  assign _0613_ = _0533_ ? 1'h0 : _0612_;
  assign _0614_ = _0534_ ? 1'h0 : _0613_;
  assign _0615_ = _0535_ ? 1'h0 : _0614_;
  assign _0616_ = _0536_ ? \u_frontend.u_npc.branch_is_call_i : _0615_;
  assign _0617_ = _0537_ ? \u_frontend.u_npc.branch_is_call_i : _0616_;
  assign _0618_ = _0538_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] ;
  assign _0619_ = _0539_ ? 1'h0 : _0618_;
  assign _0620_ = _0540_ ? 1'h0 : _0619_;
  assign _0621_ = _0541_ ? 1'h0 : _0620_;
  assign _0622_ = _0542_ ? 1'h0 : _0621_;
  assign _0623_ = _0543_ ? 1'h0 : _0622_;
  assign _0624_ = _0544_ ? 1'h0 : _0623_;
  assign _0625_ = _0545_ ? 1'h0 : _0624_;
  assign _0626_ = _0546_ ? \u_frontend.u_npc.branch_is_call_i : _0625_;
  assign _0627_ = _0547_ ? \u_frontend.u_npc.branch_is_call_i : _0626_;
  assign _0628_ = _0548_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] ;
  assign _0629_ = _0549_ ? 1'h0 : _0628_;
  assign _0630_ = _0550_ ? 1'h0 : _0629_;
  assign _0631_ = _0551_ ? 1'h0 : _0630_;
  assign _0632_ = _0552_ ? 1'h0 : _0631_;
  assign _0633_ = _0553_ ? 1'h0 : _0632_;
  assign _0634_ = _0554_ ? 1'h0 : _0633_;
  assign _0635_ = _0555_ ? 1'h0 : _0634_;
  assign _0636_ = _0556_ ? \u_frontend.u_npc.branch_is_call_i : _0635_;
  assign _0637_ = _0557_ ? \u_frontend.u_npc.branch_is_call_i : _0636_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[0] <= _0567_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[1] <= _0577_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[2] <= _0587_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[3] <= _0597_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[4] <= _0607_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[5] <= _0617_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[6] <= _0627_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_q[7] <= _0637_;
  assign _3009_ = 1'h0 ? _0639_ : _0638_;
  assign _0638_ = 1'h0 ? _0641_ : _0640_;
  assign _0639_ = 1'h0 ? _0643_ : _0642_;
  assign _0640_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0641_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0642_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0643_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3010_ = 1'h0 ? _0645_ : _0644_;
  assign _0644_ = 1'h0 ? _0647_ : _0646_;
  assign _0645_ = 1'h0 ? _0649_ : _0648_;
  assign _0646_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0647_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0648_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0649_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3011_ = 1'h0 ? _0651_ : _0650_;
  assign _0650_ = 1'h1 ? _0653_ : _0652_;
  assign _0651_ = 1'h1 ? _0655_ : _0654_;
  assign _0652_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0653_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0654_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0655_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3012_ = 1'h0 ? _0657_ : _0656_;
  assign _0656_ = 1'h1 ? _0659_ : _0658_;
  assign _0657_ = 1'h1 ? _0661_ : _0660_;
  assign _0658_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0659_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0660_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0661_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3013_ = 1'h1 ? _0663_ : _0662_;
  assign _0662_ = 1'h0 ? _0665_ : _0664_;
  assign _0663_ = 1'h0 ? _0667_ : _0666_;
  assign _0664_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0665_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0666_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0667_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3014_ = 1'h1 ? _0669_ : _0668_;
  assign _0668_ = 1'h0 ? _0671_ : _0670_;
  assign _0669_ = 1'h0 ? _0673_ : _0672_;
  assign _0670_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0671_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0672_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0673_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3015_ = 1'h1 ? _0675_ : _0674_;
  assign _0674_ = 1'h1 ? _0677_ : _0676_;
  assign _0675_ = 1'h1 ? _0679_ : _0678_;
  assign _0676_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0677_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0678_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0679_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _3016_ = 1'h1 ? _0681_ : _0680_;
  assign _0680_ = 1'h1 ? _0683_ : _0682_;
  assign _0681_ = 1'h1 ? _0685_ : _0684_;
  assign _0682_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0683_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0684_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0685_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _0686_ = _0001_ & _2827_[1];
  assign _0687_ = _0002_ & _2827_[1];
  assign _0688_ = _0004_ & _2827_[1];
  assign _0689_ = _0005_ & _2827_[1];
  assign _0690_ = _0007_ & _2827_[1];
  assign _0691_ = _0008_ & _2827_[1];
  assign _0692_ = _0010_ & _2827_[1];
  assign _0693_ = _0011_ & _2827_[1];
  assign _0694_ = _0093_ & _2832_;
  assign _0695_ = _0095_ & _2833_;
  assign _0696_ = _0014_ & _2827_[1];
  assign _0697_ = _0015_ & _2827_[1];
  assign _0698_ = _0016_ & _2827_[1];
  assign _0699_ = _0017_ & _2827_[1];
  assign _0700_ = _0018_ & _2827_[1];
  assign _0701_ = _0019_ & _2827_[1];
  assign _0702_ = _0020_ & _2827_[1];
  assign _0703_ = _0021_ & _2827_[1];
  assign _0704_ = _0096_ & _2832_;
  assign _0705_ = _0097_ & _2833_;
  assign _0706_ = _0024_ & _2827_[1];
  assign _0707_ = _0025_ & _2827_[1];
  assign _0708_ = _0027_ & _2827_[1];
  assign _0709_ = _0028_ & _2827_[1];
  assign _0710_ = _0030_ & _2827_[1];
  assign _0711_ = _0031_ & _2827_[1];
  assign _0712_ = _0033_ & _2827_[1];
  assign _0713_ = _0034_ & _2827_[1];
  assign _0714_ = _0099_ & _2832_;
  assign _0715_ = _0101_ & _2833_;
  assign _0716_ = _0037_ & _2827_[1];
  assign _0717_ = _0038_ & _2827_[1];
  assign _0718_ = _0039_ & _2827_[1];
  assign _0719_ = _0040_ & _2827_[1];
  assign _0720_ = _0041_ & _2827_[1];
  assign _0721_ = _0042_ & _2827_[1];
  assign _0722_ = _0043_ & _2827_[1];
  assign _0723_ = _0044_ & _2827_[1];
  assign _0724_ = _0102_ & _2832_;
  assign _0725_ = _0103_ & _2833_;
  assign _0726_ = _0047_ & _2827_[1];
  assign _0727_ = _0048_ & _2827_[1];
  assign _0728_ = _0050_ & _2827_[1];
  assign _0729_ = _0051_ & _2827_[1];
  assign _0730_ = _0053_ & _2827_[1];
  assign _0731_ = _0054_ & _2827_[1];
  assign _0732_ = _0056_ & _2827_[1];
  assign _0733_ = _0057_ & _2827_[1];
  assign _0734_ = _0105_ & _2832_;
  assign _0735_ = _0107_ & _2833_;
  assign _0736_ = _0060_ & _2827_[1];
  assign _0737_ = _0061_ & _2827_[1];
  assign _0738_ = _0062_ & _2827_[1];
  assign _0739_ = _0063_ & _2827_[1];
  assign _0740_ = _0064_ & _2827_[1];
  assign _0741_ = _0065_ & _2827_[1];
  assign _0742_ = _0066_ & _2827_[1];
  assign _0743_ = _0067_ & _2827_[1];
  assign _0744_ = _0108_ & _2832_;
  assign _0745_ = _0109_ & _2833_;
  assign _0746_ = _0070_ & _2827_[1];
  assign _0747_ = _0071_ & _2827_[1];
  assign _0748_ = _0073_ & _2827_[1];
  assign _0749_ = _0074_ & _2827_[1];
  assign _0750_ = _0076_ & _2827_[1];
  assign _0751_ = _0077_ & _2827_[1];
  assign _0752_ = _0079_ & _2827_[1];
  assign _0753_ = _0080_ & _2827_[1];
  assign _0754_ = _0111_ & _2832_;
  assign _0755_ = _0113_ & _2833_;
  assign _0756_ = _0083_ & _2827_[1];
  assign _0757_ = _0084_ & _2827_[1];
  assign _0758_ = _0085_ & _2827_[1];
  assign _0759_ = _0086_ & _2827_[1];
  assign _0760_ = _0087_ & _2827_[1];
  assign _0761_ = _0088_ & _2827_[1];
  assign _0762_ = _0089_ & _2827_[1];
  assign _0763_ = _0090_ & _2827_[1];
  assign _0764_ = _0114_ & _2832_;
  assign _0765_ = _0115_ & _2833_;
  assign _0766_ = _0686_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] ;
  assign _0767_ = _0687_ ? 1'h0 : _0766_;
  assign _0768_ = _0688_ ? 1'h0 : _0767_;
  assign _0769_ = _0689_ ? 1'h0 : _0768_;
  assign _0770_ = _0690_ ? 1'h0 : _0769_;
  assign _0771_ = _0691_ ? 1'h0 : _0770_;
  assign _0772_ = _0692_ ? 1'h0 : _0771_;
  assign _0773_ = _0693_ ? 1'h0 : _0772_;
  assign _0774_ = _0694_ ? \u_frontend.u_npc.branch_is_jmp_i : _0773_;
  assign _0775_ = _0695_ ? \u_frontend.u_npc.branch_is_jmp_i : _0774_;
  assign _0776_ = _0696_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] ;
  assign _0777_ = _0697_ ? 1'h0 : _0776_;
  assign _0778_ = _0698_ ? 1'h0 : _0777_;
  assign _0779_ = _0699_ ? 1'h0 : _0778_;
  assign _0780_ = _0700_ ? 1'h0 : _0779_;
  assign _0781_ = _0701_ ? 1'h0 : _0780_;
  assign _0782_ = _0702_ ? 1'h0 : _0781_;
  assign _0783_ = _0703_ ? 1'h0 : _0782_;
  assign _0784_ = _0704_ ? \u_frontend.u_npc.branch_is_jmp_i : _0783_;
  assign _0785_ = _0705_ ? \u_frontend.u_npc.branch_is_jmp_i : _0784_;
  assign _0786_ = _0706_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] ;
  assign _0787_ = _0707_ ? 1'h0 : _0786_;
  assign _0788_ = _0708_ ? 1'h0 : _0787_;
  assign _0789_ = _0709_ ? 1'h0 : _0788_;
  assign _0790_ = _0710_ ? 1'h0 : _0789_;
  assign _0791_ = _0711_ ? 1'h0 : _0790_;
  assign _0792_ = _0712_ ? 1'h0 : _0791_;
  assign _0793_ = _0713_ ? 1'h0 : _0792_;
  assign _0794_ = _0714_ ? \u_frontend.u_npc.branch_is_jmp_i : _0793_;
  assign _0795_ = _0715_ ? \u_frontend.u_npc.branch_is_jmp_i : _0794_;
  assign _0796_ = _0716_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] ;
  assign _0797_ = _0717_ ? 1'h0 : _0796_;
  assign _0798_ = _0718_ ? 1'h0 : _0797_;
  assign _0799_ = _0719_ ? 1'h0 : _0798_;
  assign _0800_ = _0720_ ? 1'h0 : _0799_;
  assign _0801_ = _0721_ ? 1'h0 : _0800_;
  assign _0802_ = _0722_ ? 1'h0 : _0801_;
  assign _0803_ = _0723_ ? 1'h0 : _0802_;
  assign _0804_ = _0724_ ? \u_frontend.u_npc.branch_is_jmp_i : _0803_;
  assign _0805_ = _0725_ ? \u_frontend.u_npc.branch_is_jmp_i : _0804_;
  assign _0806_ = _0726_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] ;
  assign _0807_ = _0727_ ? 1'h0 : _0806_;
  assign _0808_ = _0728_ ? 1'h0 : _0807_;
  assign _0809_ = _0729_ ? 1'h0 : _0808_;
  assign _0810_ = _0730_ ? 1'h0 : _0809_;
  assign _0811_ = _0731_ ? 1'h0 : _0810_;
  assign _0812_ = _0732_ ? 1'h0 : _0811_;
  assign _0813_ = _0733_ ? 1'h0 : _0812_;
  assign _0814_ = _0734_ ? \u_frontend.u_npc.branch_is_jmp_i : _0813_;
  assign _0815_ = _0735_ ? \u_frontend.u_npc.branch_is_jmp_i : _0814_;
  assign _0816_ = _0736_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] ;
  assign _0817_ = _0737_ ? 1'h0 : _0816_;
  assign _0818_ = _0738_ ? 1'h0 : _0817_;
  assign _0819_ = _0739_ ? 1'h0 : _0818_;
  assign _0820_ = _0740_ ? 1'h0 : _0819_;
  assign _0821_ = _0741_ ? 1'h0 : _0820_;
  assign _0822_ = _0742_ ? 1'h0 : _0821_;
  assign _0823_ = _0743_ ? 1'h0 : _0822_;
  assign _0824_ = _0744_ ? \u_frontend.u_npc.branch_is_jmp_i : _0823_;
  assign _0825_ = _0745_ ? \u_frontend.u_npc.branch_is_jmp_i : _0824_;
  assign _0826_ = _0746_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] ;
  assign _0827_ = _0747_ ? 1'h0 : _0826_;
  assign _0828_ = _0748_ ? 1'h0 : _0827_;
  assign _0829_ = _0749_ ? 1'h0 : _0828_;
  assign _0830_ = _0750_ ? 1'h0 : _0829_;
  assign _0831_ = _0751_ ? 1'h0 : _0830_;
  assign _0832_ = _0752_ ? 1'h0 : _0831_;
  assign _0833_ = _0753_ ? 1'h0 : _0832_;
  assign _0834_ = _0754_ ? \u_frontend.u_npc.branch_is_jmp_i : _0833_;
  assign _0835_ = _0755_ ? \u_frontend.u_npc.branch_is_jmp_i : _0834_;
  assign _0836_ = _0756_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] ;
  assign _0837_ = _0757_ ? 1'h0 : _0836_;
  assign _0838_ = _0758_ ? 1'h0 : _0837_;
  assign _0839_ = _0759_ ? 1'h0 : _0838_;
  assign _0840_ = _0760_ ? 1'h0 : _0839_;
  assign _0841_ = _0761_ ? 1'h0 : _0840_;
  assign _0842_ = _0762_ ? 1'h0 : _0841_;
  assign _0843_ = _0763_ ? 1'h0 : _0842_;
  assign _0844_ = _0764_ ? \u_frontend.u_npc.branch_is_jmp_i : _0843_;
  assign _0845_ = _0765_ ? \u_frontend.u_npc.branch_is_jmp_i : _0844_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[0] <= _0775_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[1] <= _0785_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[2] <= _0795_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[3] <= _0805_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[4] <= _0815_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[5] <= _0825_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[6] <= _0835_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_q[7] <= _0845_;
  assign _3017_ = 1'h0 ? _0847_ : _0846_;
  assign _0846_ = 1'h0 ? _0849_ : _0848_;
  assign _0847_ = 1'h0 ? _0851_ : _0850_;
  assign _0848_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0849_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0850_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0851_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3018_ = 1'h0 ? _0853_ : _0852_;
  assign _0852_ = 1'h0 ? _0855_ : _0854_;
  assign _0853_ = 1'h0 ? _0857_ : _0856_;
  assign _0854_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0855_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0856_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0857_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3019_ = 1'h0 ? _0859_ : _0858_;
  assign _0858_ = 1'h1 ? _0861_ : _0860_;
  assign _0859_ = 1'h1 ? _0863_ : _0862_;
  assign _0860_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0861_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0862_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0863_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3020_ = 1'h0 ? _0865_ : _0864_;
  assign _0864_ = 1'h1 ? _0867_ : _0866_;
  assign _0865_ = 1'h1 ? _0869_ : _0868_;
  assign _0866_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0867_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0868_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0869_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3021_ = 1'h1 ? _0871_ : _0870_;
  assign _0870_ = 1'h0 ? _0873_ : _0872_;
  assign _0871_ = 1'h0 ? _0875_ : _0874_;
  assign _0872_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0873_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0874_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0875_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3022_ = 1'h1 ? _0877_ : _0876_;
  assign _0876_ = 1'h0 ? _0879_ : _0878_;
  assign _0877_ = 1'h0 ? _0881_ : _0880_;
  assign _0878_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0879_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0880_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0881_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3023_ = 1'h1 ? _0883_ : _0882_;
  assign _0882_ = 1'h1 ? _0885_ : _0884_;
  assign _0883_ = 1'h1 ? _0887_ : _0886_;
  assign _0884_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0885_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0886_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0887_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _3024_ = 1'h1 ? _0889_ : _0888_;
  assign _0888_ = 1'h1 ? _0891_ : _0890_;
  assign _0889_ = 1'h1 ? _0893_ : _0892_;
  assign _0890_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0891_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0892_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _0893_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _0894_ = _0001_ & _2827_[1];
  assign _0895_ = _0002_ & _2827_[1];
  assign _0896_ = _0004_ & _2827_[1];
  assign _0897_ = _0005_ & _2827_[1];
  assign _0898_ = _0007_ & _2827_[1];
  assign _0899_ = _0008_ & _2827_[1];
  assign _0900_ = _0010_ & _2827_[1];
  assign _0901_ = _0011_ & _2827_[1];
  assign _0902_ = _0093_ & _2832_;
  assign _0903_ = _0095_ & _2833_;
  assign _0904_ = _0014_ & _2827_[1];
  assign _0905_ = _0015_ & _2827_[1];
  assign _0906_ = _0016_ & _2827_[1];
  assign _0907_ = _0017_ & _2827_[1];
  assign _0908_ = _0018_ & _2827_[1];
  assign _0909_ = _0019_ & _2827_[1];
  assign _0910_ = _0020_ & _2827_[1];
  assign _0911_ = _0021_ & _2827_[1];
  assign _0912_ = _0096_ & _2832_;
  assign _0913_ = _0097_ & _2833_;
  assign _0914_ = _0024_ & _2827_[1];
  assign _0915_ = _0025_ & _2827_[1];
  assign _0916_ = _0027_ & _2827_[1];
  assign _0917_ = _0028_ & _2827_[1];
  assign _0918_ = _0030_ & _2827_[1];
  assign _0919_ = _0031_ & _2827_[1];
  assign _0920_ = _0033_ & _2827_[1];
  assign _0921_ = _0034_ & _2827_[1];
  assign _0922_ = _0099_ & _2832_;
  assign _0923_ = _0101_ & _2833_;
  assign _0924_ = _0037_ & _2827_[1];
  assign _0925_ = _0038_ & _2827_[1];
  assign _0926_ = _0039_ & _2827_[1];
  assign _0927_ = _0040_ & _2827_[1];
  assign _0928_ = _0041_ & _2827_[1];
  assign _0929_ = _0042_ & _2827_[1];
  assign _0930_ = _0043_ & _2827_[1];
  assign _0931_ = _0044_ & _2827_[1];
  assign _0932_ = _0102_ & _2832_;
  assign _0933_ = _0103_ & _2833_;
  assign _0934_ = _0047_ & _2827_[1];
  assign _0935_ = _0048_ & _2827_[1];
  assign _0936_ = _0050_ & _2827_[1];
  assign _0937_ = _0051_ & _2827_[1];
  assign _0938_ = _0053_ & _2827_[1];
  assign _0939_ = _0054_ & _2827_[1];
  assign _0940_ = _0056_ & _2827_[1];
  assign _0941_ = _0057_ & _2827_[1];
  assign _0942_ = _0105_ & _2832_;
  assign _0943_ = _0107_ & _2833_;
  assign _0944_ = _0060_ & _2827_[1];
  assign _0945_ = _0061_ & _2827_[1];
  assign _0946_ = _0062_ & _2827_[1];
  assign _0947_ = _0063_ & _2827_[1];
  assign _0948_ = _0064_ & _2827_[1];
  assign _0949_ = _0065_ & _2827_[1];
  assign _0950_ = _0066_ & _2827_[1];
  assign _0951_ = _0067_ & _2827_[1];
  assign _0952_ = _0108_ & _2832_;
  assign _0953_ = _0109_ & _2833_;
  assign _0954_ = _0070_ & _2827_[1];
  assign _0955_ = _0071_ & _2827_[1];
  assign _0956_ = _0073_ & _2827_[1];
  assign _0957_ = _0074_ & _2827_[1];
  assign _0958_ = _0076_ & _2827_[1];
  assign _0959_ = _0077_ & _2827_[1];
  assign _0960_ = _0079_ & _2827_[1];
  assign _0961_ = _0080_ & _2827_[1];
  assign _0962_ = _0111_ & _2832_;
  assign _0963_ = _0113_ & _2833_;
  assign _0964_ = _0083_ & _2827_[1];
  assign _0965_ = _0084_ & _2827_[1];
  assign _0966_ = _0085_ & _2827_[1];
  assign _0967_ = _0086_ & _2827_[1];
  assign _0968_ = _0087_ & _2827_[1];
  assign _0969_ = _0088_ & _2827_[1];
  assign _0970_ = _0089_ & _2827_[1];
  assign _0971_ = _0090_ & _2827_[1];
  assign _0972_ = _0114_ & _2832_;
  assign _0973_ = _0115_ & _2833_;
  assign _0974_ = _0894_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] ;
  assign _0975_ = _0895_ ? 1'h0 : _0974_;
  assign _0976_ = _0896_ ? 1'h0 : _0975_;
  assign _0977_ = _0897_ ? 1'h0 : _0976_;
  assign _0978_ = _0898_ ? 1'h0 : _0977_;
  assign _0979_ = _0899_ ? 1'h0 : _0978_;
  assign _0980_ = _0900_ ? 1'h0 : _0979_;
  assign _0981_ = _0901_ ? 1'h0 : _0980_;
  assign _0982_ = _0902_ ? \u_frontend.u_npc.branch_is_ret_i : _0981_;
  assign _0983_ = _0903_ ? \u_frontend.u_npc.branch_is_ret_i : _0982_;
  assign _0984_ = _0904_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] ;
  assign _0985_ = _0905_ ? 1'h0 : _0984_;
  assign _0986_ = _0906_ ? 1'h0 : _0985_;
  assign _0987_ = _0907_ ? 1'h0 : _0986_;
  assign _0988_ = _0908_ ? 1'h0 : _0987_;
  assign _0989_ = _0909_ ? 1'h0 : _0988_;
  assign _0990_ = _0910_ ? 1'h0 : _0989_;
  assign _0991_ = _0911_ ? 1'h0 : _0990_;
  assign _0992_ = _0912_ ? \u_frontend.u_npc.branch_is_ret_i : _0991_;
  assign _0993_ = _0913_ ? \u_frontend.u_npc.branch_is_ret_i : _0992_;
  assign _0994_ = _0914_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] ;
  assign _0995_ = _0915_ ? 1'h0 : _0994_;
  assign _0996_ = _0916_ ? 1'h0 : _0995_;
  assign _0997_ = _0917_ ? 1'h0 : _0996_;
  assign _0998_ = _0918_ ? 1'h0 : _0997_;
  assign _0999_ = _0919_ ? 1'h0 : _0998_;
  assign _1000_ = _0920_ ? 1'h0 : _0999_;
  assign _1001_ = _0921_ ? 1'h0 : _1000_;
  assign _1002_ = _0922_ ? \u_frontend.u_npc.branch_is_ret_i : _1001_;
  assign _1003_ = _0923_ ? \u_frontend.u_npc.branch_is_ret_i : _1002_;
  assign _1004_ = _0924_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] ;
  assign _1005_ = _0925_ ? 1'h0 : _1004_;
  assign _1006_ = _0926_ ? 1'h0 : _1005_;
  assign _1007_ = _0927_ ? 1'h0 : _1006_;
  assign _1008_ = _0928_ ? 1'h0 : _1007_;
  assign _1009_ = _0929_ ? 1'h0 : _1008_;
  assign _1010_ = _0930_ ? 1'h0 : _1009_;
  assign _1011_ = _0931_ ? 1'h0 : _1010_;
  assign _1012_ = _0932_ ? \u_frontend.u_npc.branch_is_ret_i : _1011_;
  assign _1013_ = _0933_ ? \u_frontend.u_npc.branch_is_ret_i : _1012_;
  assign _1014_ = _0934_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] ;
  assign _1015_ = _0935_ ? 1'h0 : _1014_;
  assign _1016_ = _0936_ ? 1'h0 : _1015_;
  assign _1017_ = _0937_ ? 1'h0 : _1016_;
  assign _1018_ = _0938_ ? 1'h0 : _1017_;
  assign _1019_ = _0939_ ? 1'h0 : _1018_;
  assign _1020_ = _0940_ ? 1'h0 : _1019_;
  assign _1021_ = _0941_ ? 1'h0 : _1020_;
  assign _1022_ = _0942_ ? \u_frontend.u_npc.branch_is_ret_i : _1021_;
  assign _1023_ = _0943_ ? \u_frontend.u_npc.branch_is_ret_i : _1022_;
  assign _1024_ = _0944_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] ;
  assign _1025_ = _0945_ ? 1'h0 : _1024_;
  assign _1026_ = _0946_ ? 1'h0 : _1025_;
  assign _1027_ = _0947_ ? 1'h0 : _1026_;
  assign _1028_ = _0948_ ? 1'h0 : _1027_;
  assign _1029_ = _0949_ ? 1'h0 : _1028_;
  assign _1030_ = _0950_ ? 1'h0 : _1029_;
  assign _1031_ = _0951_ ? 1'h0 : _1030_;
  assign _1032_ = _0952_ ? \u_frontend.u_npc.branch_is_ret_i : _1031_;
  assign _1033_ = _0953_ ? \u_frontend.u_npc.branch_is_ret_i : _1032_;
  assign _1034_ = _0954_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] ;
  assign _1035_ = _0955_ ? 1'h0 : _1034_;
  assign _1036_ = _0956_ ? 1'h0 : _1035_;
  assign _1037_ = _0957_ ? 1'h0 : _1036_;
  assign _1038_ = _0958_ ? 1'h0 : _1037_;
  assign _1039_ = _0959_ ? 1'h0 : _1038_;
  assign _1040_ = _0960_ ? 1'h0 : _1039_;
  assign _1041_ = _0961_ ? 1'h0 : _1040_;
  assign _1042_ = _0962_ ? \u_frontend.u_npc.branch_is_ret_i : _1041_;
  assign _1043_ = _0963_ ? \u_frontend.u_npc.branch_is_ret_i : _1042_;
  assign _1044_ = _0964_ ? 1'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] ;
  assign _1045_ = _0965_ ? 1'h0 : _1044_;
  assign _1046_ = _0966_ ? 1'h0 : _1045_;
  assign _1047_ = _0967_ ? 1'h0 : _1046_;
  assign _1048_ = _0968_ ? 1'h0 : _1047_;
  assign _1049_ = _0969_ ? 1'h0 : _1048_;
  assign _1050_ = _0970_ ? 1'h0 : _1049_;
  assign _1051_ = _0971_ ? 1'h0 : _1050_;
  assign _1052_ = _0972_ ? \u_frontend.u_npc.branch_is_ret_i : _1051_;
  assign _1053_ = _0973_ ? \u_frontend.u_npc.branch_is_ret_i : _1052_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[0] <= _0983_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[1] <= _0993_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[2] <= _1003_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[3] <= _1013_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[4] <= _1023_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[5] <= _1033_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[6] <= _1043_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_q[7] <= _1053_;
  assign _3025_ = 1'h0 ? _1055_ : _1054_;
  assign _1054_ = 1'h0 ? _1057_ : _1056_;
  assign _1055_ = 1'h0 ? _1059_ : _1058_;
  assign _1056_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1057_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1058_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1059_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3026_ = 1'h0 ? _1061_ : _1060_;
  assign _1060_ = 1'h0 ? _1063_ : _1062_;
  assign _1061_ = 1'h0 ? _1065_ : _1064_;
  assign _1062_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1063_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1064_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1065_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3027_ = 1'h0 ? _1067_ : _1066_;
  assign _1066_ = 1'h1 ? _1069_ : _1068_;
  assign _1067_ = 1'h1 ? _1071_ : _1070_;
  assign _1068_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1069_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1070_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1071_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3028_ = 1'h0 ? _1073_ : _1072_;
  assign _1072_ = 1'h1 ? _1075_ : _1074_;
  assign _1073_ = 1'h1 ? _1077_ : _1076_;
  assign _1074_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1075_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1076_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1077_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3029_ = 1'h1 ? _1079_ : _1078_;
  assign _1078_ = 1'h0 ? _1081_ : _1080_;
  assign _1079_ = 1'h0 ? _1083_ : _1082_;
  assign _1080_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1081_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1082_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1083_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3030_ = 1'h1 ? _1085_ : _1084_;
  assign _1084_ = 1'h0 ? _1087_ : _1086_;
  assign _1085_ = 1'h0 ? _1089_ : _1088_;
  assign _1086_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1087_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1088_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1089_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3031_ = 1'h1 ? _1091_ : _1090_;
  assign _1090_ = 1'h1 ? _1093_ : _1092_;
  assign _1091_ = 1'h1 ? _1095_ : _1094_;
  assign _1092_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1093_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1094_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1095_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _3032_ = 1'h1 ? _1097_ : _1096_;
  assign _1096_ = 1'h1 ? _1099_ : _1098_;
  assign _1097_ = 1'h1 ? _1101_ : _1100_;
  assign _1098_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1099_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1100_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1101_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _1102_ = _0001_ & _2827_[1];
  assign _1103_ = _0002_ & _2827_[1];
  assign _1104_ = _0004_ & _2827_[1];
  assign _1105_ = _0005_ & _2827_[1];
  assign _1106_ = _0007_ & _2827_[1];
  assign _1107_ = _0008_ & _2827_[1];
  assign _1108_ = _0010_ & _2827_[1];
  assign _1109_ = _0011_ & _2827_[1];
  assign _1110_ = _0093_ & _2832_;
  assign _1111_ = _0095_ & _2833_;
  assign _1112_ = _0014_ & _2827_[1];
  assign _1113_ = _0015_ & _2827_[1];
  assign _1114_ = _0016_ & _2827_[1];
  assign _1115_ = _0017_ & _2827_[1];
  assign _1116_ = _0018_ & _2827_[1];
  assign _1117_ = _0019_ & _2827_[1];
  assign _1118_ = _0020_ & _2827_[1];
  assign _1119_ = _0021_ & _2827_[1];
  assign _1120_ = _0096_ & _2832_;
  assign _1121_ = _0097_ & _2833_;
  assign _1122_ = _0024_ & _2827_[1];
  assign _1123_ = _0025_ & _2827_[1];
  assign _1124_ = _0027_ & _2827_[1];
  assign _1125_ = _0028_ & _2827_[1];
  assign _1126_ = _0030_ & _2827_[1];
  assign _1127_ = _0031_ & _2827_[1];
  assign _1128_ = _0033_ & _2827_[1];
  assign _1129_ = _0034_ & _2827_[1];
  assign _1130_ = _0099_ & _2832_;
  assign _1131_ = _0101_ & _2833_;
  assign _1132_ = _0037_ & _2827_[1];
  assign _1133_ = _0038_ & _2827_[1];
  assign _1134_ = _0039_ & _2827_[1];
  assign _1135_ = _0040_ & _2827_[1];
  assign _1136_ = _0041_ & _2827_[1];
  assign _1137_ = _0042_ & _2827_[1];
  assign _1138_ = _0043_ & _2827_[1];
  assign _1139_ = _0044_ & _2827_[1];
  assign _1140_ = _0102_ & _2832_;
  assign _1141_ = _0103_ & _2833_;
  assign _1142_ = _0047_ & _2827_[1];
  assign _1143_ = _0048_ & _2827_[1];
  assign _1144_ = _0050_ & _2827_[1];
  assign _1145_ = _0051_ & _2827_[1];
  assign _1146_ = _0053_ & _2827_[1];
  assign _1147_ = _0054_ & _2827_[1];
  assign _1148_ = _0056_ & _2827_[1];
  assign _1149_ = _0057_ & _2827_[1];
  assign _1150_ = _0105_ & _2832_;
  assign _1151_ = _0107_ & _2833_;
  assign _1152_ = _0060_ & _2827_[1];
  assign _1153_ = _0061_ & _2827_[1];
  assign _1154_ = _0062_ & _2827_[1];
  assign _1155_ = _0063_ & _2827_[1];
  assign _1156_ = _0064_ & _2827_[1];
  assign _1157_ = _0065_ & _2827_[1];
  assign _1158_ = _0066_ & _2827_[1];
  assign _1159_ = _0067_ & _2827_[1];
  assign _1160_ = _0108_ & _2832_;
  assign _1161_ = _0109_ & _2833_;
  assign _1162_ = _0070_ & _2827_[1];
  assign _1163_ = _0071_ & _2827_[1];
  assign _1164_ = _0073_ & _2827_[1];
  assign _1165_ = _0074_ & _2827_[1];
  assign _1166_ = _0076_ & _2827_[1];
  assign _1167_ = _0077_ & _2827_[1];
  assign _1168_ = _0079_ & _2827_[1];
  assign _1169_ = _0080_ & _2827_[1];
  assign _1170_ = _0111_ & _2832_;
  assign _1171_ = _0113_ & _2833_;
  assign _1172_ = _0083_ & _2827_[1];
  assign _1173_ = _0084_ & _2827_[1];
  assign _1174_ = _0085_ & _2827_[1];
  assign _1175_ = _0086_ & _2827_[1];
  assign _1176_ = _0087_ & _2827_[1];
  assign _1177_ = _0088_ & _2827_[1];
  assign _1178_ = _0089_ & _2827_[1];
  assign _1179_ = _0090_ & _2827_[1];
  assign _1180_ = _0114_ & _2832_;
  assign _1181_ = _0115_ & _2833_;
  assign _1182_ = _1102_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] ;
  assign _1183_ = _1103_ ? 32'h00000000 : _1182_;
  assign _1184_ = _1104_ ? 32'h00000000 : _1183_;
  assign _1185_ = _1105_ ? 32'h00000000 : _1184_;
  assign _1186_ = _1106_ ? 32'h00000000 : _1185_;
  assign _1187_ = _1107_ ? 32'h00000000 : _1186_;
  assign _1188_ = _1108_ ? 32'h00000000 : _1187_;
  assign _1189_ = _1109_ ? 32'h00000000 : _1188_;
  assign _1190_ = _1110_ ? \u_frontend.u_npc.branch_source_i : _1189_;
  assign _1191_ = _1111_ ? \u_frontend.u_npc.branch_source_i : _1190_;
  assign _1192_ = _1112_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] ;
  assign _1193_ = _1113_ ? 32'h00000000 : _1192_;
  assign _1194_ = _1114_ ? 32'h00000000 : _1193_;
  assign _1195_ = _1115_ ? 32'h00000000 : _1194_;
  assign _1196_ = _1116_ ? 32'h00000000 : _1195_;
  assign _1197_ = _1117_ ? 32'h00000000 : _1196_;
  assign _1198_ = _1118_ ? 32'h00000000 : _1197_;
  assign _1199_ = _1119_ ? 32'h00000000 : _1198_;
  assign _1200_ = _1120_ ? \u_frontend.u_npc.branch_source_i : _1199_;
  assign _1201_ = _1121_ ? \u_frontend.u_npc.branch_source_i : _1200_;
  assign _1202_ = _1122_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] ;
  assign _1203_ = _1123_ ? 32'h00000000 : _1202_;
  assign _1204_ = _1124_ ? 32'h00000000 : _1203_;
  assign _1205_ = _1125_ ? 32'h00000000 : _1204_;
  assign _1206_ = _1126_ ? 32'h00000000 : _1205_;
  assign _1207_ = _1127_ ? 32'h00000000 : _1206_;
  assign _1208_ = _1128_ ? 32'h00000000 : _1207_;
  assign _1209_ = _1129_ ? 32'h00000000 : _1208_;
  assign _1210_ = _1130_ ? \u_frontend.u_npc.branch_source_i : _1209_;
  assign _1211_ = _1131_ ? \u_frontend.u_npc.branch_source_i : _1210_;
  assign _1212_ = _1132_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] ;
  assign _1213_ = _1133_ ? 32'h00000000 : _1212_;
  assign _1214_ = _1134_ ? 32'h00000000 : _1213_;
  assign _1215_ = _1135_ ? 32'h00000000 : _1214_;
  assign _1216_ = _1136_ ? 32'h00000000 : _1215_;
  assign _1217_ = _1137_ ? 32'h00000000 : _1216_;
  assign _1218_ = _1138_ ? 32'h00000000 : _1217_;
  assign _1219_ = _1139_ ? 32'h00000000 : _1218_;
  assign _1220_ = _1140_ ? \u_frontend.u_npc.branch_source_i : _1219_;
  assign _1221_ = _1141_ ? \u_frontend.u_npc.branch_source_i : _1220_;
  assign _1222_ = _1142_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] ;
  assign _1223_ = _1143_ ? 32'h00000000 : _1222_;
  assign _1224_ = _1144_ ? 32'h00000000 : _1223_;
  assign _1225_ = _1145_ ? 32'h00000000 : _1224_;
  assign _1226_ = _1146_ ? 32'h00000000 : _1225_;
  assign _1227_ = _1147_ ? 32'h00000000 : _1226_;
  assign _1228_ = _1148_ ? 32'h00000000 : _1227_;
  assign _1229_ = _1149_ ? 32'h00000000 : _1228_;
  assign _1230_ = _1150_ ? \u_frontend.u_npc.branch_source_i : _1229_;
  assign _1231_ = _1151_ ? \u_frontend.u_npc.branch_source_i : _1230_;
  assign _1232_ = _1152_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] ;
  assign _1233_ = _1153_ ? 32'h00000000 : _1232_;
  assign _1234_ = _1154_ ? 32'h00000000 : _1233_;
  assign _1235_ = _1155_ ? 32'h00000000 : _1234_;
  assign _1236_ = _1156_ ? 32'h00000000 : _1235_;
  assign _1237_ = _1157_ ? 32'h00000000 : _1236_;
  assign _1238_ = _1158_ ? 32'h00000000 : _1237_;
  assign _1239_ = _1159_ ? 32'h00000000 : _1238_;
  assign _1240_ = _1160_ ? \u_frontend.u_npc.branch_source_i : _1239_;
  assign _1241_ = _1161_ ? \u_frontend.u_npc.branch_source_i : _1240_;
  assign _1242_ = _1162_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] ;
  assign _1243_ = _1163_ ? 32'h00000000 : _1242_;
  assign _1244_ = _1164_ ? 32'h00000000 : _1243_;
  assign _1245_ = _1165_ ? 32'h00000000 : _1244_;
  assign _1246_ = _1166_ ? 32'h00000000 : _1245_;
  assign _1247_ = _1167_ ? 32'h00000000 : _1246_;
  assign _1248_ = _1168_ ? 32'h00000000 : _1247_;
  assign _1249_ = _1169_ ? 32'h00000000 : _1248_;
  assign _1250_ = _1170_ ? \u_frontend.u_npc.branch_source_i : _1249_;
  assign _1251_ = _1171_ ? \u_frontend.u_npc.branch_source_i : _1250_;
  assign _1252_ = _1172_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] ;
  assign _1253_ = _1173_ ? 32'h00000000 : _1252_;
  assign _1254_ = _1174_ ? 32'h00000000 : _1253_;
  assign _1255_ = _1175_ ? 32'h00000000 : _1254_;
  assign _1256_ = _1176_ ? 32'h00000000 : _1255_;
  assign _1257_ = _1177_ ? 32'h00000000 : _1256_;
  assign _1258_ = _1178_ ? 32'h00000000 : _1257_;
  assign _1259_ = _1179_ ? 32'h00000000 : _1258_;
  assign _1260_ = _1180_ ? \u_frontend.u_npc.branch_source_i : _1259_;
  assign _1261_ = _1181_ ? \u_frontend.u_npc.branch_source_i : _1260_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[0] <= _1191_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[1] <= _1201_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[2] <= _1211_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[3] <= _1221_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[4] <= _1231_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[5] <= _1241_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[6] <= _1251_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_pc_q[7] <= _1261_;
  assign _3033_ = 1'h0 ? _1263_ : _1262_;
  assign _1262_ = 1'h0 ? _1265_ : _1264_;
  assign _1263_ = 1'h0 ? _1267_ : _1266_;
  assign _1264_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1265_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1266_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1267_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3034_ = 1'h0 ? _1269_ : _1268_;
  assign _1268_ = 1'h0 ? _1271_ : _1270_;
  assign _1269_ = 1'h0 ? _1273_ : _1272_;
  assign _1270_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1271_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1272_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1273_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3035_ = 1'h0 ? _1275_ : _1274_;
  assign _1274_ = 1'h1 ? _1277_ : _1276_;
  assign _1275_ = 1'h1 ? _1279_ : _1278_;
  assign _1276_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1277_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1278_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1279_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3036_ = 1'h0 ? _1281_ : _1280_;
  assign _1280_ = 1'h1 ? _1283_ : _1282_;
  assign _1281_ = 1'h1 ? _1285_ : _1284_;
  assign _1282_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1283_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1284_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1285_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3037_ = 1'h1 ? _1287_ : _1286_;
  assign _1286_ = 1'h0 ? _1289_ : _1288_;
  assign _1287_ = 1'h0 ? _1291_ : _1290_;
  assign _1288_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1289_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1290_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1291_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3038_ = 1'h1 ? _1293_ : _1292_;
  assign _1292_ = 1'h0 ? _1295_ : _1294_;
  assign _1293_ = 1'h0 ? _1297_ : _1296_;
  assign _1294_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1295_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1296_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1297_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3039_ = 1'h1 ? _1299_ : _1298_;
  assign _1298_ = 1'h1 ? _1301_ : _1300_;
  assign _1299_ = 1'h1 ? _1303_ : _1302_;
  assign _1300_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1301_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1302_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1303_ = 1'h0 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _3040_ = 1'h1 ? _1305_ : _1304_;
  assign _1304_ = 1'h1 ? _1307_ : _1306_;
  assign _1305_ = 1'h1 ? _1309_ : _1308_;
  assign _1306_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1307_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1308_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1309_ = 1'h1 ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _1310_ = _0001_ & _2827_[1];
  assign _1311_ = _0002_ & _2827_[1];
  assign _1312_ = _0004_ & _2827_[1];
  assign _1313_ = _0005_ & _2827_[1];
  assign _1314_ = _0007_ & _2827_[1];
  assign _1315_ = _0008_ & _2827_[1];
  assign _1316_ = _0010_ & _2827_[1];
  assign _1317_ = _0011_ & _2827_[1];
  assign _1318_ = _0093_ & _2834_[31];
  assign _1319_ = _0095_ & _2833_;
  assign _1320_ = _0014_ & _2827_[1];
  assign _1321_ = _0015_ & _2827_[1];
  assign _1322_ = _0016_ & _2827_[1];
  assign _1323_ = _0017_ & _2827_[1];
  assign _1324_ = _0018_ & _2827_[1];
  assign _1325_ = _0019_ & _2827_[1];
  assign _1326_ = _0020_ & _2827_[1];
  assign _1327_ = _0021_ & _2827_[1];
  assign _1328_ = _0096_ & _2834_[31];
  assign _1329_ = _0097_ & _2833_;
  assign _1330_ = _0024_ & _2827_[1];
  assign _1331_ = _0025_ & _2827_[1];
  assign _1332_ = _0027_ & _2827_[1];
  assign _1333_ = _0028_ & _2827_[1];
  assign _1334_ = _0030_ & _2827_[1];
  assign _1335_ = _0031_ & _2827_[1];
  assign _1336_ = _0033_ & _2827_[1];
  assign _1337_ = _0034_ & _2827_[1];
  assign _1338_ = _0099_ & _2834_[31];
  assign _1339_ = _0101_ & _2833_;
  assign _1340_ = _0037_ & _2827_[1];
  assign _1341_ = _0038_ & _2827_[1];
  assign _1342_ = _0039_ & _2827_[1];
  assign _1343_ = _0040_ & _2827_[1];
  assign _1344_ = _0041_ & _2827_[1];
  assign _1345_ = _0042_ & _2827_[1];
  assign _1346_ = _0043_ & _2827_[1];
  assign _1347_ = _0044_ & _2827_[1];
  assign _1348_ = _0102_ & _2834_[31];
  assign _1349_ = _0103_ & _2833_;
  assign _1350_ = _0047_ & _2827_[1];
  assign _1351_ = _0048_ & _2827_[1];
  assign _1352_ = _0050_ & _2827_[1];
  assign _1353_ = _0051_ & _2827_[1];
  assign _1354_ = _0053_ & _2827_[1];
  assign _1355_ = _0054_ & _2827_[1];
  assign _1356_ = _0056_ & _2827_[1];
  assign _1357_ = _0057_ & _2827_[1];
  assign _1358_ = _0105_ & _2834_[31];
  assign _1359_ = _0107_ & _2833_;
  assign _1360_ = _0060_ & _2827_[1];
  assign _1361_ = _0061_ & _2827_[1];
  assign _1362_ = _0062_ & _2827_[1];
  assign _1363_ = _0063_ & _2827_[1];
  assign _1364_ = _0064_ & _2827_[1];
  assign _1365_ = _0065_ & _2827_[1];
  assign _1366_ = _0066_ & _2827_[1];
  assign _1367_ = _0067_ & _2827_[1];
  assign _1368_ = _0108_ & _2834_[31];
  assign _1369_ = _0109_ & _2833_;
  assign _1370_ = _0070_ & _2827_[1];
  assign _1371_ = _0071_ & _2827_[1];
  assign _1372_ = _0073_ & _2827_[1];
  assign _1373_ = _0074_ & _2827_[1];
  assign _1374_ = _0076_ & _2827_[1];
  assign _1375_ = _0077_ & _2827_[1];
  assign _1376_ = _0079_ & _2827_[1];
  assign _1377_ = _0080_ & _2827_[1];
  assign _1378_ = _0111_ & _2834_[31];
  assign _1379_ = _0113_ & _2833_;
  assign _1380_ = _0083_ & _2827_[1];
  assign _1381_ = _0084_ & _2827_[1];
  assign _1382_ = _0085_ & _2827_[1];
  assign _1383_ = _0086_ & _2827_[1];
  assign _1384_ = _0087_ & _2827_[1];
  assign _1385_ = _0088_ & _2827_[1];
  assign _1386_ = _0089_ & _2827_[1];
  assign _1387_ = _0090_ & _2827_[1];
  assign _1388_ = _0114_ & _2834_[31];
  assign _1389_ = _0115_ & _2833_;
  assign _1390_ = _1310_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] ;
  assign _1391_ = _1311_ ? 32'h00000000 : _1390_;
  assign _1392_ = _1312_ ? 32'h00000000 : _1391_;
  assign _1393_ = _1313_ ? 32'h00000000 : _1392_;
  assign _1394_ = _1314_ ? 32'h00000000 : _1393_;
  assign _1395_ = _1315_ ? 32'h00000000 : _1394_;
  assign _1396_ = _1316_ ? 32'h00000000 : _1395_;
  assign _1397_ = _1317_ ? 32'h00000000 : _1396_;
  assign _1398_ = _1318_ ? \u_frontend.u_npc.branch_pc_i : _1397_;
  assign _1399_ = _1319_ ? \u_frontend.u_npc.branch_pc_i : _1398_;
  assign _1400_ = _1320_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] ;
  assign _1401_ = _1321_ ? 32'h00000000 : _1400_;
  assign _1402_ = _1322_ ? 32'h00000000 : _1401_;
  assign _1403_ = _1323_ ? 32'h00000000 : _1402_;
  assign _1404_ = _1324_ ? 32'h00000000 : _1403_;
  assign _1405_ = _1325_ ? 32'h00000000 : _1404_;
  assign _1406_ = _1326_ ? 32'h00000000 : _1405_;
  assign _1407_ = _1327_ ? 32'h00000000 : _1406_;
  assign _1408_ = _1328_ ? \u_frontend.u_npc.branch_pc_i : _1407_;
  assign _1409_ = _1329_ ? \u_frontend.u_npc.branch_pc_i : _1408_;
  assign _1410_ = _1330_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] ;
  assign _1411_ = _1331_ ? 32'h00000000 : _1410_;
  assign _1412_ = _1332_ ? 32'h00000000 : _1411_;
  assign _1413_ = _1333_ ? 32'h00000000 : _1412_;
  assign _1414_ = _1334_ ? 32'h00000000 : _1413_;
  assign _1415_ = _1335_ ? 32'h00000000 : _1414_;
  assign _1416_ = _1336_ ? 32'h00000000 : _1415_;
  assign _1417_ = _1337_ ? 32'h00000000 : _1416_;
  assign _1418_ = _1338_ ? \u_frontend.u_npc.branch_pc_i : _1417_;
  assign _1419_ = _1339_ ? \u_frontend.u_npc.branch_pc_i : _1418_;
  assign _1420_ = _1340_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] ;
  assign _1421_ = _1341_ ? 32'h00000000 : _1420_;
  assign _1422_ = _1342_ ? 32'h00000000 : _1421_;
  assign _1423_ = _1343_ ? 32'h00000000 : _1422_;
  assign _1424_ = _1344_ ? 32'h00000000 : _1423_;
  assign _1425_ = _1345_ ? 32'h00000000 : _1424_;
  assign _1426_ = _1346_ ? 32'h00000000 : _1425_;
  assign _1427_ = _1347_ ? 32'h00000000 : _1426_;
  assign _1428_ = _1348_ ? \u_frontend.u_npc.branch_pc_i : _1427_;
  assign _1429_ = _1349_ ? \u_frontend.u_npc.branch_pc_i : _1428_;
  assign _1430_ = _1350_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] ;
  assign _1431_ = _1351_ ? 32'h00000000 : _1430_;
  assign _1432_ = _1352_ ? 32'h00000000 : _1431_;
  assign _1433_ = _1353_ ? 32'h00000000 : _1432_;
  assign _1434_ = _1354_ ? 32'h00000000 : _1433_;
  assign _1435_ = _1355_ ? 32'h00000000 : _1434_;
  assign _1436_ = _1356_ ? 32'h00000000 : _1435_;
  assign _1437_ = _1357_ ? 32'h00000000 : _1436_;
  assign _1438_ = _1358_ ? \u_frontend.u_npc.branch_pc_i : _1437_;
  assign _1439_ = _1359_ ? \u_frontend.u_npc.branch_pc_i : _1438_;
  assign _1440_ = _1360_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] ;
  assign _1441_ = _1361_ ? 32'h00000000 : _1440_;
  assign _1442_ = _1362_ ? 32'h00000000 : _1441_;
  assign _1443_ = _1363_ ? 32'h00000000 : _1442_;
  assign _1444_ = _1364_ ? 32'h00000000 : _1443_;
  assign _1445_ = _1365_ ? 32'h00000000 : _1444_;
  assign _1446_ = _1366_ ? 32'h00000000 : _1445_;
  assign _1447_ = _1367_ ? 32'h00000000 : _1446_;
  assign _1448_ = _1368_ ? \u_frontend.u_npc.branch_pc_i : _1447_;
  assign _1449_ = _1369_ ? \u_frontend.u_npc.branch_pc_i : _1448_;
  assign _1450_ = _1370_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] ;
  assign _1451_ = _1371_ ? 32'h00000000 : _1450_;
  assign _1452_ = _1372_ ? 32'h00000000 : _1451_;
  assign _1453_ = _1373_ ? 32'h00000000 : _1452_;
  assign _1454_ = _1374_ ? 32'h00000000 : _1453_;
  assign _1455_ = _1375_ ? 32'h00000000 : _1454_;
  assign _1456_ = _1376_ ? 32'h00000000 : _1455_;
  assign _1457_ = _1377_ ? 32'h00000000 : _1456_;
  assign _1458_ = _1378_ ? \u_frontend.u_npc.branch_pc_i : _1457_;
  assign _1459_ = _1379_ ? \u_frontend.u_npc.branch_pc_i : _1458_;
  assign _1460_ = _1380_ ? 32'h00000000 : \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] ;
  assign _1461_ = _1381_ ? 32'h00000000 : _1460_;
  assign _1462_ = _1382_ ? 32'h00000000 : _1461_;
  assign _1463_ = _1383_ ? 32'h00000000 : _1462_;
  assign _1464_ = _1384_ ? 32'h00000000 : _1463_;
  assign _1465_ = _1385_ ? 32'h00000000 : _1464_;
  assign _1466_ = _1386_ ? 32'h00000000 : _1465_;
  assign _1467_ = _1387_ ? 32'h00000000 : _1466_;
  assign _1468_ = _1388_ ? \u_frontend.u_npc.branch_pc_i : _1467_;
  assign _1469_ = _1389_ ? \u_frontend.u_npc.branch_pc_i : _1468_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[0] <= _1399_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[1] <= _1409_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[2] <= _1419_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[3] <= _1429_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[4] <= _1439_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[5] <= _1449_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[6] <= _1459_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.btb_target_q[7] <= _1469_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.ras_pc_pred_w = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [2] ? _1471_ : _1470_;
  assign _1470_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [1] ? _1473_ : _1472_;
  assign _1471_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [1] ? _1475_ : _1474_;
  assign _1472_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [0] ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[1] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[0] ;
  assign _1473_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [0] ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[3] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[2] ;
  assign _1474_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [0] ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[5] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[4] ;
  assign _1475_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q [0] ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[7] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[6] ;
  assign _1476_ = _0001_ & _2827_[1];
  assign _1477_ = _0002_ & _2827_[1];
  assign _1478_ = _0004_ & _2827_[1];
  assign _1479_ = _0005_ & _2827_[1];
  assign _1480_ = _0007_ & _2827_[1];
  assign _1481_ = _0008_ & _2827_[1];
  assign _1482_ = _0010_ & _2827_[1];
  assign _1483_ = _0011_ & _2827_[1];
  assign _1484_ = _0117_ & _2836_[31];
  assign _1485_ = _0117_ & _2838_[31];
  assign _1486_ = _0014_ & _2827_[1];
  assign _1487_ = _0015_ & _2827_[1];
  assign _1488_ = _0016_ & _2827_[1];
  assign _1489_ = _0017_ & _2827_[1];
  assign _1490_ = _0018_ & _2827_[1];
  assign _1491_ = _0019_ & _2827_[1];
  assign _1492_ = _0020_ & _2827_[1];
  assign _1493_ = _0021_ & _2827_[1];
  assign _1494_ = _0118_ & _2836_[31];
  assign _1495_ = _0118_ & _2838_[31];
  assign _1496_ = _0024_ & _2827_[1];
  assign _1497_ = _0025_ & _2827_[1];
  assign _1498_ = _0027_ & _2827_[1];
  assign _1499_ = _0028_ & _2827_[1];
  assign _1500_ = _0030_ & _2827_[1];
  assign _1501_ = _0031_ & _2827_[1];
  assign _1502_ = _0033_ & _2827_[1];
  assign _1503_ = _0034_ & _2827_[1];
  assign _1504_ = _0120_ & _2836_[31];
  assign _1505_ = _0120_ & _2838_[31];
  assign _1506_ = _0037_ & _2827_[1];
  assign _1507_ = _0038_ & _2827_[1];
  assign _1508_ = _0039_ & _2827_[1];
  assign _1509_ = _0040_ & _2827_[1];
  assign _1510_ = _0041_ & _2827_[1];
  assign _1511_ = _0042_ & _2827_[1];
  assign _1512_ = _0043_ & _2827_[1];
  assign _1513_ = _0044_ & _2827_[1];
  assign _1514_ = _0121_ & _2836_[31];
  assign _1515_ = _0121_ & _2838_[31];
  assign _1516_ = _0047_ & _2827_[1];
  assign _1517_ = _0048_ & _2827_[1];
  assign _1518_ = _0050_ & _2827_[1];
  assign _1519_ = _0051_ & _2827_[1];
  assign _1520_ = _0053_ & _2827_[1];
  assign _1521_ = _0054_ & _2827_[1];
  assign _1522_ = _0056_ & _2827_[1];
  assign _1523_ = _0057_ & _2827_[1];
  assign _1524_ = _0123_ & _2836_[31];
  assign _1525_ = _0123_ & _2838_[31];
  assign _1526_ = _0060_ & _2827_[1];
  assign _1527_ = _0061_ & _2827_[1];
  assign _1528_ = _0062_ & _2827_[1];
  assign _1529_ = _0063_ & _2827_[1];
  assign _1530_ = _0064_ & _2827_[1];
  assign _1531_ = _0065_ & _2827_[1];
  assign _1532_ = _0066_ & _2827_[1];
  assign _1533_ = _0067_ & _2827_[1];
  assign _1534_ = _0124_ & _2836_[31];
  assign _1535_ = _0124_ & _2838_[31];
  assign _1536_ = _0070_ & _2827_[1];
  assign _1537_ = _0071_ & _2827_[1];
  assign _1538_ = _0073_ & _2827_[1];
  assign _1539_ = _0074_ & _2827_[1];
  assign _1540_ = _0076_ & _2827_[1];
  assign _1541_ = _0077_ & _2827_[1];
  assign _1542_ = _0079_ & _2827_[1];
  assign _1543_ = _0080_ & _2827_[1];
  assign _1544_ = _0126_ & _2836_[31];
  assign _1545_ = _0126_ & _2838_[31];
  assign _1546_ = _0083_ & _2827_[1];
  assign _1547_ = _0084_ & _2827_[1];
  assign _1548_ = _0085_ & _2827_[1];
  assign _1549_ = _0086_ & _2827_[1];
  assign _1550_ = _0087_ & _2827_[1];
  assign _1551_ = _0088_ & _2827_[1];
  assign _1552_ = _0089_ & _2827_[1];
  assign _1553_ = _0090_ & _2827_[1];
  assign _1554_ = _0127_ & _2836_[31];
  assign _1555_ = _0127_ & _2838_[31];
  assign _1556_ = _1476_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[0] ;
  assign _1557_ = _1477_ ? 32'h00000001 : _1556_;
  assign _1558_ = _1478_ ? 32'h00000001 : _1557_;
  assign _1559_ = _1479_ ? 32'h00000001 : _1558_;
  assign _1560_ = _1480_ ? 32'h00000001 : _1559_;
  assign _1561_ = _1481_ ? 32'h00000001 : _1560_;
  assign _1562_ = _1482_ ? 32'h00000001 : _1561_;
  assign _1563_ = _1483_ ? 32'h00000001 : _1562_;
  assign _1564_ = _1484_ ? _2835_ : _1563_;
  assign _1565_ = _1485_ ? _2837_ : _1564_;
  assign _1566_ = _1486_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[1] ;
  assign _1567_ = _1487_ ? 32'h00000001 : _1566_;
  assign _1568_ = _1488_ ? 32'h00000001 : _1567_;
  assign _1569_ = _1489_ ? 32'h00000001 : _1568_;
  assign _1570_ = _1490_ ? 32'h00000001 : _1569_;
  assign _1571_ = _1491_ ? 32'h00000001 : _1570_;
  assign _1572_ = _1492_ ? 32'h00000001 : _1571_;
  assign _1573_ = _1493_ ? 32'h00000001 : _1572_;
  assign _1574_ = _1494_ ? _2835_ : _1573_;
  assign _1575_ = _1495_ ? _2837_ : _1574_;
  assign _1576_ = _1496_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[2] ;
  assign _1577_ = _1497_ ? 32'h00000001 : _1576_;
  assign _1578_ = _1498_ ? 32'h00000001 : _1577_;
  assign _1579_ = _1499_ ? 32'h00000001 : _1578_;
  assign _1580_ = _1500_ ? 32'h00000001 : _1579_;
  assign _1581_ = _1501_ ? 32'h00000001 : _1580_;
  assign _1582_ = _1502_ ? 32'h00000001 : _1581_;
  assign _1583_ = _1503_ ? 32'h00000001 : _1582_;
  assign _1584_ = _1504_ ? _2835_ : _1583_;
  assign _1585_ = _1505_ ? _2837_ : _1584_;
  assign _1586_ = _1506_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[3] ;
  assign _1587_ = _1507_ ? 32'h00000001 : _1586_;
  assign _1588_ = _1508_ ? 32'h00000001 : _1587_;
  assign _1589_ = _1509_ ? 32'h00000001 : _1588_;
  assign _1590_ = _1510_ ? 32'h00000001 : _1589_;
  assign _1591_ = _1511_ ? 32'h00000001 : _1590_;
  assign _1592_ = _1512_ ? 32'h00000001 : _1591_;
  assign _1593_ = _1513_ ? 32'h00000001 : _1592_;
  assign _1594_ = _1514_ ? _2835_ : _1593_;
  assign _1595_ = _1515_ ? _2837_ : _1594_;
  assign _1596_ = _1516_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[4] ;
  assign _1597_ = _1517_ ? 32'h00000001 : _1596_;
  assign _1598_ = _1518_ ? 32'h00000001 : _1597_;
  assign _1599_ = _1519_ ? 32'h00000001 : _1598_;
  assign _1600_ = _1520_ ? 32'h00000001 : _1599_;
  assign _1601_ = _1521_ ? 32'h00000001 : _1600_;
  assign _1602_ = _1522_ ? 32'h00000001 : _1601_;
  assign _1603_ = _1523_ ? 32'h00000001 : _1602_;
  assign _1604_ = _1524_ ? _2835_ : _1603_;
  assign _1605_ = _1525_ ? _2837_ : _1604_;
  assign _1606_ = _1526_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[5] ;
  assign _1607_ = _1527_ ? 32'h00000001 : _1606_;
  assign _1608_ = _1528_ ? 32'h00000001 : _1607_;
  assign _1609_ = _1529_ ? 32'h00000001 : _1608_;
  assign _1610_ = _1530_ ? 32'h00000001 : _1609_;
  assign _1611_ = _1531_ ? 32'h00000001 : _1610_;
  assign _1612_ = _1532_ ? 32'h00000001 : _1611_;
  assign _1613_ = _1533_ ? 32'h00000001 : _1612_;
  assign _1614_ = _1534_ ? _2835_ : _1613_;
  assign _1615_ = _1535_ ? _2837_ : _1614_;
  assign _1616_ = _1536_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[6] ;
  assign _1617_ = _1537_ ? 32'h00000001 : _1616_;
  assign _1618_ = _1538_ ? 32'h00000001 : _1617_;
  assign _1619_ = _1539_ ? 32'h00000001 : _1618_;
  assign _1620_ = _1540_ ? 32'h00000001 : _1619_;
  assign _1621_ = _1541_ ? 32'h00000001 : _1620_;
  assign _1622_ = _1542_ ? 32'h00000001 : _1621_;
  assign _1623_ = _1543_ ? 32'h00000001 : _1622_;
  assign _1624_ = _1544_ ? _2835_ : _1623_;
  assign _1625_ = _1545_ ? _2837_ : _1624_;
  assign _1626_ = _1546_ ? 32'h00000001 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[7] ;
  assign _1627_ = _1547_ ? 32'h00000001 : _1626_;
  assign _1628_ = _1548_ ? 32'h00000001 : _1627_;
  assign _1629_ = _1549_ ? 32'h00000001 : _1628_;
  assign _1630_ = _1550_ ? 32'h00000001 : _1629_;
  assign _1631_ = _1551_ ? 32'h00000001 : _1630_;
  assign _1632_ = _1552_ ? 32'h00000001 : _1631_;
  assign _1633_ = _1553_ ? 32'h00000001 : _1632_;
  assign _1634_ = _1554_ ? _2835_ : _1633_;
  assign _1635_ = _1555_ ? _2837_ : _1634_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[0] <= _1565_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[1] <= _1575_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[2] <= _1585_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[3] <= _1595_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[4] <= _1605_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[5] <= _1615_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[6] <= _1625_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_stack_q[7] <= _1635_;
  assign \u_lsu.u_lsu_request.data_out_o = \u_lsu.u_lsu_request.rd_ptr_q ? \u_lsu.u_lsu_request.ram_q[1] : \u_lsu.u_lsu_request.ram_q[0] ;
  assign _1636_ = _0128_ & _4130_[35];
  assign _1637_ = _0129_ & _4130_[35];
  assign _1638_ = _0160_ & _4131_[35];
  assign _1639_ = _0131_ & _4130_[35];
  assign _1640_ = _0132_ & _4130_[35];
  assign _1641_ = _0161_ & _4131_[35];
  assign _1642_ = _1636_ ? 36'h000000000 : \u_lsu.u_lsu_request.ram_q[0] ;
  assign _1643_ = _1637_ ? 36'h000000000 : _1642_;
  logic [35:0] fangyuan6;
  assign fangyuan6 = { \u_lsu.mem_addr_q , \u_lsu.mem_ls_q , \u_lsu.mem_xh_q , \u_lsu.mem_xb_q , \u_lsu.mem_load_q };
  assign _1644_ = _1638_ ? fangyuan6 : _1643_;
  assign _1645_ = _1639_ ? 36'h000000000 : \u_lsu.u_lsu_request.ram_q[1] ;
  assign _1646_ = _1640_ ? 36'h000000000 : _1645_;
  logic [35:0] fangyuan7;
  assign fangyuan7 = { \u_lsu.mem_addr_q , \u_lsu.mem_ls_q , \u_lsu.mem_xh_q , \u_lsu.mem_xb_q , \u_lsu.mem_load_q };
  assign _1647_ = _1641_ ? fangyuan7 : _1646_;
  always @(posedge clk_i)
      \u_lsu.u_lsu_request.ram_q[0] <= _1644_;
  always @(posedge clk_i)
      \u_lsu.u_lsu_request.ram_q[1] <= _1647_;
  assign _1657_ = 5'h18 + \u_csr.u_csrfile.csr_mpriv_q ;
  assign _1658_ = \u_csr.opcode_opcode_i & 15'h707f;
  assign _1659_ = \u_csr.opcode_opcode_i & 32'hffffffff;
  assign _1660_ = \u_csr.opcode_opcode_i & 32'hdfffffff;
  assign _1661_ = \u_csr.csr_rdata_w & _1683_;
  assign _1662_ = _1708_ & _1684_;
  assign _1663_ = \u_csr.opcode_opcode_i & 32'hfe007fff;
  assign _1664_ = _1658_ == 13'h100f;
  assign _1665_ = \u_csr.opcode_opcode_i [31:20] == 9'h180;
  assign _1666_ = _1659_ == 7'h73;
  assign _1667_ = _1660_ == 29'h10200073;
  assign _1668_ = _1659_ == 21'h100073;
  assign _1669_ = _1658_ == 13'h1073;
  assign _1670_ = _1658_ == 14'h2073;
  assign _1671_ = _1658_ == 14'h3073;
  assign _1672_ = _1658_ == 15'h5073;
  assign _1673_ = _1658_ == 15'h6073;
  assign _1674_ = _1658_ == 15'h7073;
  assign _1675_ = _1663_ == 29'h12000073;
  assign \u_csr.ifence_w = \u_csr.opcode_valid_i && _1664_;
  assign _1676_ = \u_csr.opcode_valid_i && _1678_;
  assign _1677_ = _1676_ && \u_csr.csr_write_r ;
  assign \u_csr.satp_update_w = _1677_ && _1665_;
  assign _1679_ = \u_csr.set_r && \u_csr.clr_r ;
  assign \u_csr.csrrw_w = \u_csr.opcode_valid_i && _1669_;
  assign \u_csr.csrrs_w = \u_csr.opcode_valid_i && _1670_;
  assign \u_csr.csrrc_w = \u_csr.opcode_valid_i && _1671_;
  assign \u_csr.csrrwi_w = \u_csr.opcode_valid_i && _1672_;
  assign \u_csr.csrrsi_w = \u_csr.opcode_valid_i && _1673_;
  assign \u_csr.csrrci_w = \u_csr.opcode_valid_i && _1674_;
  assign \u_csr.sfence_w = \u_csr.opcode_valid_i && _1675_;
  assign _1678_ = \u_csr.set_r || \u_csr.clr_r ;
  assign _1680_ = \u_csr.satp_update_w || \u_csr.ifence_w ;
  assign _1681_ = _1680_ || \u_csr.sfence_w ;
  assign _1682_ = | \u_csr.opcode_opcode_i [19:15];
  assign _1683_ = ~ \u_csr.data_r ;
  assign _1684_ = ~ \u_csr.interrupt_inhibit_i ;
  assign _1685_ = \u_csr.csrrw_w | \u_csr.csrrs_w ;
  assign _1686_ = _1685_ | \u_csr.csrrwi_w ;
  assign \u_csr.set_r = _1686_ | \u_csr.csrrsi_w ;
  assign _1687_ = \u_csr.csrrw_w | \u_csr.csrrc_w ;
  assign _1688_ = _1687_ | \u_csr.csrrwi_w ;
  assign \u_csr.clr_r = _1688_ | \u_csr.csrrci_w ;
  assign _1689_ = _1682_ | \u_csr.csrrw_w ;
  assign \u_csr.csr_write_r = _1689_ | \u_csr.csrrwi_w ;
  assign _1690_ = \u_csr.csrrwi_w | \u_csr.csrrsi_w ;
  assign _1691_ = _1690_ | \u_csr.csrrci_w ;
  assign _1692_ = \u_csr.csr_rdata_w | \u_csr.data_r ;
  always @(posedge clk_i)
      \u_csr.branch_q <= _1648_;
  always @(posedge clk_i)
      \u_csr.branch_target_q <= _1649_;
  always @(posedge clk_i)
      \u_csr.reset_q <= _1655_;
  always @(posedge clk_i)
      \u_csr.ifence_q <= _1652_;
  always @(posedge clk_i)
      \u_csr.take_interrupt_q <= _1656_;
  always @(posedge clk_i)
      \u_csr.rd_valid_e1_q <= _1654_;
  always @(posedge clk_i)
      \u_csr.rd_result_e1_q <= _1653_;
  always @(posedge clk_i)
      \u_csr.csr_wdata_e1_q <= _1650_;
  always @(posedge clk_i)
      \u_csr.exception_e1_q <= _1651_;
  assign _1655_ = rst_i ? 1'h1 : 1'h0;
  assign _1693_ = \u_csr.reset_q ? reset_vector_i : \u_csr.csr_target_w ;
  assign _1649_ = rst_i ? 32'h00000000 : _1693_;
  assign _1694_ = \u_csr.reset_q ? 1'h1 : \u_csr.csr_branch_w ;
  assign _1648_ = rst_i ? 1'h0 : _1694_;
  assign _1652_ = rst_i ? 1'h0 : \u_csr.ifence_w ;
  assign _1656_ = rst_i ? 1'h0 : _1662_;
  assign _1695_ = _1681_ ? 6'h31 : 6'h00;
  assign _1696_ = \u_csr.opcode_invalid_i ? 6'h12 : _1695_;
  assign _1697_ = _1668_ ? 6'h13 : _1696_;
  assign _1698_ = _1667_ ? 6'h30 : _1697_;
  assign _1699_ = _1666_ ? _1657_ : _1698_;
  assign _1700_ = \u_csr.opcode_valid_i ? _1699_ : 6'h00;
  assign _1651_ = rst_i ? 6'h00 : _1700_;
  assign _1701_ = \u_csr.clr_r ? _1661_ : \u_csr.csr_wdata_e1_q ;
  assign _1702_ = \u_csr.set_r ? _1692_ : _1701_;
  assign _1703_ = _1679_ ? \u_csr.data_r : _1702_;
  assign _1704_ = \u_csr.opcode_valid_i ? _1703_ : 32'h00000000;
  assign _1650_ = rst_i ? 32'h00000000 : _1704_;
  assign _1705_ = \u_csr.opcode_invalid_i ? \u_csr.opcode_opcode_i : \u_csr.csr_rdata_w ;
  assign _1706_ = \u_csr.opcode_valid_i ? _1705_ : 32'h00000000;
  assign _1653_ = rst_i ? 32'h00000000 : _1706_;
  assign _1707_ = \u_csr.opcode_valid_i ? _1678_ : 1'h0;
  assign _1654_ = rst_i ? 1'h0 : _1707_;
  logic [31:0] fangyuan8;
  assign fangyuan8 = { \u_csr.interrupt_w [0], \u_csr.interrupt_w [1], \u_csr.interrupt_w [2], \u_csr.interrupt_w [3], \u_csr.interrupt_w [4], \u_csr.interrupt_w [5], \u_csr.interrupt_w [6], \u_csr.interrupt_w [7], \u_csr.interrupt_w [8], \u_csr.interrupt_w [9], \u_csr.interrupt_w [10], \u_csr.interrupt_w [11], \u_csr.interrupt_w [12], \u_csr.interrupt_w [13], \u_csr.interrupt_w [14], \u_csr.interrupt_w [15], \u_csr.interrupt_w [16], \u_csr.interrupt_w [17], \u_csr.interrupt_w [18], \u_csr.interrupt_w [19], \u_csr.interrupt_w [20], \u_csr.interrupt_w [21], \u_csr.interrupt_w [22], \u_csr.interrupt_w [23], \u_csr.interrupt_w [24], \u_csr.interrupt_w [25], \u_csr.interrupt_w [26], \u_csr.interrupt_w [27], \u_csr.interrupt_w [28], \u_csr.interrupt_w [29], \u_csr.interrupt_w [30], \u_csr.interrupt_w [31] };
  assign _1708_ = | fangyuan8;
  logic [31:0] fangyuan9;
  assign fangyuan9 = { 27'h0000000, \u_csr.opcode_opcode_i [19:15] };
  assign \u_csr.data_r = _1691_ ? fangyuan9 : \u_csr.opcode_ra_operand_i ;
  assign \u_csr.u_csrfile.csr_waddr_i = \u_issue.u_pipe0_ctrl.csr_wr_wb_q ? \u_issue.u_pipe0_ctrl.opcode_wb_q [31:20] : 12'h000;
  assign \u_csr.u_csrfile.csr_mcycle_r = \u_csr.u_csrfile.csr_mcycle_q + 1'h1;
  assign _1774_ = \u_csr.u_csrfile.exception_pc_i + 3'h4;
  assign \u_csr.u_csrfile.irq_pending_r = \u_csr.u_csrfile.csr_mip_q & \u_csr.u_csrfile.csr_mie_q ;
  assign _1775_ = \u_csr.u_csrfile.csr_mscratch_q & 32'hffffffff;
  assign _1776_ = \u_csr.u_csrfile.csr_mepc_q & 32'hffffffff;
  assign _1777_ = \u_csr.u_csrfile.csr_mtvec_q & 32'hffffffff;
  assign _1778_ = \u_csr.u_csrfile.csr_mcause_q & 32'h8000000f;
  assign _1779_ = \u_csr.u_csrfile.csr_mtval_q & 32'hffffffff;
  assign _1780_ = \u_csr.u_csrfile.csr_sr_q & 32'hffffffff;
  assign _1781_ = \u_csr.u_csrfile.csr_mip_q & 12'haaa;
  assign _1782_ = \u_csr.u_csrfile.csr_mie_q & 12'haaa;
  assign _1783_ = \u_csr.u_csrfile.exception_i & 6'h30;
  assign _1784_ = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q & 32'hffffffff;
  assign _1785_ = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q & 32'h8000000f;
  assign _1786_ = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q & 12'haaa;
  assign _1787_ = \u_csr.u_csrfile.csr_sr_q & 32'hfffbfecc;
  assign _1788_ = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q & 19'h40133;
  assign _1789_ = \u_csr.u_csrfile.csr_mip_q & 32'hfffffddd;
  assign _1790_ = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q & 10'h222;
  assign _1791_ = \u_csr.u_csrfile.csr_mie_q & 32'hfffffddd;
  assign _1792_ = \u_csr.opcode_opcode_i [31:20] == 10'h344;
  assign _1793_ = \u_csr.opcode_opcode_i [31:20] == 9'h144;
  assign _1794_ = \u_csr.u_csrfile.csr_waddr_i == 10'h344;
  assign _1795_ = \u_csr.u_csrfile.csr_waddr_i == 9'h144;
  assign \u_csr.u_csrfile.is_exception_w = _1783_ == 5'h10;
  assign _1796_ = _1783_ == 6'h20;
  assign _1797_ = \u_csr.u_csrfile.irq_priv_q == 2'h3;
  assign _1798_ = \u_csr.u_csrfile.csr_mpriv_q == 1'h1;
  assign _1799_ = \u_csr.u_csrfile.exception_i == 6'h30;
  assign _1800_ = \u_csr.u_csrfile.csr_mpriv_q == 2'h3;
  assign _1801_ = \u_csr.u_csrfile.csr_mcycle_q == \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign _1802_ = \u_csr.u_csrfile.exception_i == 6'h20;
  assign _1803_ = \u_csr.u_csrfile.exception_i == 6'h31;
  assign _1804_ = \u_csr.opcode_valid_i && _1792_;
  assign _1805_ = \u_csr.opcode_valid_i && _1793_;
  assign _1806_ = intr_i && \u_csr.u_csrfile.csr_mtimecmp_q [11];
  assign _1807_ = intr_i && _1814_;
  assign _1808_ = 1'h0 && \u_csr.u_csrfile.csr_mtimecmp_q [7];
  assign _1809_ = 1'h0 && _1815_;
  assign _1810_ = $signed(32'h00000000) && _1801_;
  assign _1811_ = _1804_ || _1805_;
  assign _1812_ = _1794_ || _1795_;
  assign _1813_ = _1812_ || _1848_;
  assign _1814_ = ~ \u_csr.u_csrfile.csr_mtimecmp_q [11];
  assign _1815_ = ~ \u_csr.u_csrfile.csr_mtimecmp_q [7];
  assign _1816_ = _1804_ | _1805_;
  assign \u_csr.u_csrfile.buffer_mip_w = _1816_ | \u_csr.u_csrfile.csr_mip_upd_q ;
  assign _1817_ = _1787_ | _1788_;
  assign _1818_ = _1789_ | _1790_;
  assign _1819_ = _1791_ | _1790_;
  logic [31:0] fangyuan10;
  assign fangyuan10 = { \u_csr.u_csrfile.csr_mip_next_q [31:12], \u_csr.u_csrfile.csr_mip_next_r [11], \u_csr.u_csrfile.csr_mip_next_q [10], \u_csr.u_csrfile.csr_mip_next_r [9], \u_csr.u_csrfile.csr_mip_next_q [8], \u_csr.u_csrfile.csr_mip_next_r [7], \u_csr.u_csrfile.csr_mip_next_q [6], \u_csr.u_csrfile.csr_mip_next_r [5], \u_csr.u_csrfile.csr_mip_next_q [4:0] };
  assign \u_csr.u_csrfile.csr_mip_r = _1726_ | fangyuan10;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mepc_q <= _1711_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mcause_q <= _1709_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_sr_q <= _1719_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mtvec_q <= _1718_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mip_q <= _1714_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mie_q <= _1712_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mpriv_q <= 2'h3;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mcycle_q <= _1710_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mscratch_q <= _1716_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mtval_q <= _1717_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mtimecmp_q <= 32'h00000000;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mtime_ie_q <= 1'h0;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mip_next_q <= _1713_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.csr_mip_upd_q <= _1715_;
  always @(posedge clk_i)
      \u_csr.u_csrfile.irq_priv_q <= _1720_;
  assign _1761_ = _1803_ ? _1774_ : 32'h00000000;
  assign _1760_ = _1803_ ? 1'h1 : 1'h0;
  assign _1748_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mtvec_q : _1761_;
  assign _1747_ = \u_csr.u_csrfile.is_exception_w ? 1'h1 : _1760_;
  assign _1737_ = _1800_ ? \u_csr.u_csrfile.csr_mepc_q : \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign _1728_ = _1799_ ? _1737_ : _1748_;
  assign _1727_ = _1799_ ? 1'h1 : _1747_;
  assign \u_csr.csr_target_w = _1802_ ? _1850_ : _1728_;
  assign \u_csr.csr_branch_w = _1802_ ? 1'h1 : _1727_;
  assign _1713_ = rst_i ? 32'h00000000 : _1849_;
  assign _1717_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mtval_r ;
  assign _1716_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mscratch_r ;
  assign _1710_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mcycle_r ;
  assign _1712_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mie_r ;
  assign _1714_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mip_r ;
  assign _1718_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mtvec_r ;
  assign _1719_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_sr_r ;
  assign _1709_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mcause_r ;
  assign _1711_ = rst_i ? 32'h00000000 : \u_csr.u_csrfile.csr_mepc_r ;
  assign _1767_ = \u_csr.u_csrfile.csr_mtimecmp_q [7] ? \u_csr.u_csrfile.csr_mtime_ie_q : _1741_;
  assign _1770_ = \u_csr.u_csrfile.csr_mtimecmp_q [7] ? _1751_ : \u_csr.u_csrfile.csr_mtime_ie_q ;
  assign \u_csr.u_csrfile.csr_mip_next_r [7] = _1810_ ? _1770_ : _1751_;
  assign \u_csr.u_csrfile.csr_mip_next_r [5] = _1810_ ? _1767_ : _1741_;
  assign _1751_ = _1809_ ? 1'h1 : \u_csr.u_csrfile.csr_mip_next_q [7];
  assign _1741_ = _1808_ ? 1'h1 : \u_csr.u_csrfile.csr_mip_next_q [5];
  assign \u_csr.u_csrfile.csr_mip_next_r [11] = _1807_ ? 1'h1 : \u_csr.u_csrfile.csr_mip_next_q [11];
  assign \u_csr.u_csrfile.csr_mip_next_r [9] = _1806_ ? 1'h1 : \u_csr.u_csrfile.csr_mip_next_q [9];
  assign _1757_ = _1820_ ? _1784_ : \u_csr.u_csrfile.csr_mscratch_q ;
  assign _1820_ = \u_csr.u_csrfile.csr_waddr_i == 10'h340;
  logic [63:0] fangyuan11;
  assign fangyuan11 = { _1786_, _1819_ };
  logic [1:0] fangyuan12;
  assign fangyuan12 = { _1822_, _1821_ };
  always @(\u_csr.u_csrfile.csr_mie_q or fangyuan11 or fangyuan12) begin
    casez (fangyuan12)
      2'b?1 :
        _1755_ = fangyuan11 [31:0] ;
      2'b1? :
        _1755_ = fangyuan11 [63:32] ;
      default:
        _1755_ = \u_csr.u_csrfile.csr_mie_q ;
    endcase
  end
  assign _1821_ = \u_csr.u_csrfile.csr_waddr_i == 9'h104;
  assign _1822_ = \u_csr.u_csrfile.csr_waddr_i == 10'h304;
  logic [63:0] fangyuan13;
  assign fangyuan13 = { _1786_, _1818_ };
  logic [1:0] fangyuan14;
  assign fangyuan14 = { _1794_, _1795_ };
  always @(\u_csr.u_csrfile.csr_mip_q or fangyuan13 or fangyuan14) begin
    casez (fangyuan14)
      2'b?1 :
        _1756_ = fangyuan13 [31:0] ;
      2'b1? :
        _1756_ = fangyuan13 [63:32] ;
      default:
        _1756_ = \u_csr.u_csrfile.csr_mip_q ;
    endcase
  end
  assign _1758_ = _1823_ ? _1784_ : \u_csr.u_csrfile.csr_mtvec_q ;
  assign _1823_ = \u_csr.u_csrfile.csr_waddr_i == 10'h305;
  logic [63:0] fangyuan15;
  assign fangyuan15 = { _1784_, _1817_ };
  logic [1:0] fangyuan16;
  assign fangyuan16 = { _1825_, _1824_ };
  always @(\u_csr.u_csrfile.csr_sr_q or fangyuan15 or fangyuan16) begin
    casez (fangyuan16)
      2'b?1 :
        _1725_ = fangyuan15 [31:0] ;
      2'b1? :
        _1725_ = fangyuan15 [63:32] ;
      default:
        _1725_ = \u_csr.u_csrfile.csr_sr_q ;
    endcase
  end
  assign _1824_ = \u_csr.u_csrfile.csr_waddr_i == 9'h100;
  assign _1825_ = \u_csr.u_csrfile.csr_waddr_i == 10'h300;
  assign _1768_ = _1826_ ? _1784_ : \u_csr.u_csrfile.csr_mtval_q ;
  assign _1826_ = \u_csr.u_csrfile.csr_waddr_i == 10'h343;
  assign _1772_ = _1827_ ? _1785_ : \u_csr.u_csrfile.csr_mcause_q ;
  assign _1827_ = \u_csr.u_csrfile.csr_waddr_i == 10'h342;
  assign _1763_ = _1828_ ? _1784_ : \u_csr.u_csrfile.csr_mepc_q ;
  assign _1828_ = \u_csr.u_csrfile.csr_waddr_i == 10'h341;
  assign _1724_[31:13] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_sr_q [31:13] : _1725_[31:13];
  assign _1724_[10:8] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_sr_q [10:8] : _1725_[10:8];
  assign _1724_[6:4] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_sr_q [6:4] : _1725_[6:4];
  assign _1724_[2:0] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_sr_q [2:0] : _1725_[2:0];
  logic [31:0] fangyuan17;
  assign fangyuan17 = { 28'h0000000, \u_csr.u_csrfile.exception_i [3:0] };
  assign _1766_ = \u_csr.u_csrfile.is_exception_w ? fangyuan17 : _1772_;
  assign _1752_ = \u_csr.u_csrfile.is_exception_w ? _1764_ : _1768_;
  assign _1750_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.exception_pc_i : _1763_;
  assign _1724_[3] = \u_csr.u_csrfile.is_exception_w ? 1'h0 : _1725_[3];
  assign _1724_[12:11] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mpriv_q : _1725_[12:11];
  assign _1724_[7] = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_sr_q [3] : _1725_[7];
  assign _1743_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mscratch_q : _1757_;
  assign _1740_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mie_q : _1755_;
  assign _1742_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mip_q : _1756_;
  assign _1745_ = \u_csr.u_csrfile.is_exception_w ? \u_csr.u_csrfile.csr_mtvec_q : _1758_;
  logic [63:0] fangyuan18;
  assign fangyuan18 = { \u_csr.u_csrfile.exception_pc_i , \u_csr.u_csrfile.exception_addr_i };
  logic [1:0] fangyuan19;
  assign fangyuan19 = { _1832_, _1830_ };
  always @(32'h00000000 or fangyuan18 or fangyuan19) begin
    casez (fangyuan19)
      2'b?1 :
        _1764_ = fangyuan18 [31:0] ;
      2'b1? :
        _1764_ = fangyuan18 [63:32] ;
      default:
        _1764_ = 32'h00000000 ;
    endcase
  end
  logic [6:0] fangyuan20;
  assign fangyuan20 = { _1829_[0], _1829_[1], _1829_[2], _1829_[3], _1829_[4], _1829_[5], _1829_[6] };
  assign _1830_ = | fangyuan20;
  assign _1829_[0] = \u_csr.u_csrfile.exception_i == 5'h12;
  assign _1829_[1] = \u_csr.u_csrfile.exception_i == 5'h14;
  assign _1829_[2] = \u_csr.u_csrfile.exception_i == 5'h15;
  assign _1829_[3] = \u_csr.u_csrfile.exception_i == 5'h16;
  assign _1829_[4] = \u_csr.u_csrfile.exception_i == 5'h17;
  assign _1829_[5] = \u_csr.u_csrfile.exception_i == 5'h1d;
  assign _1829_[6] = \u_csr.u_csrfile.exception_i == 5'h1f;
  logic [2:0] fangyuan21;
  assign fangyuan21 = { _1831_[0], _1831_[1], _1831_[2] };
  assign _1832_ = | fangyuan21;
  assign _1831_[0] = \u_csr.u_csrfile.exception_i == 5'h10;
  assign _1831_[1] = \u_csr.u_csrfile.exception_i == 5'h11;
  assign _1831_[2] = \u_csr.u_csrfile.exception_i == 5'h1c;
  assign _1769_[31:13] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [31:13] : _1724_[31:13];
  assign _1769_[10:9] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [10:9] : _1724_[10:9];
  assign _1769_[6] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [6] : _1724_[6];
  assign _1769_[4] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [4] : _1724_[4];
  assign _1769_[2] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [2] : _1724_[2];
  assign _1769_[0] = _1799_ ? \u_csr.u_csrfile.csr_sr_q [0] : _1724_[0];
  assign _1722_[0] = _1800_ ? 1'h1 : \u_csr.u_csrfile.csr_sr_q [7];
  assign _1773_ = _1800_ ? \u_csr.u_csrfile.csr_sr_q [7] : \u_csr.u_csrfile.csr_sr_q [3];
  assign _1722_[1] = _1800_ ? \u_csr.u_csrfile.csr_sr_q [8] : 1'h0;
  assign _1721_ = _1800_ ? \u_csr.u_csrfile.csr_sr_q [5] : 1'h1;
  assign _1771_ = _1800_ ? \u_csr.u_csrfile.csr_sr_q [1] : \u_csr.u_csrfile.csr_sr_q [5];
  assign _1769_[12:11] = _1799_ ? _1723_ : _1724_[12:11];
  assign _1769_[8:7] = _1799_ ? _1722_ : _1724_[8:7];
  assign _1769_[5] = _1799_ ? _1721_ : _1724_[5];
  assign _1769_[3] = _1799_ ? _1773_ : _1724_[3];
  assign _1769_[1] = _1799_ ? _1771_ : _1724_[1];
  assign _1733_ = _1799_ ? \u_csr.u_csrfile.csr_mscratch_q : _1743_;
  assign _1731_ = _1799_ ? \u_csr.u_csrfile.csr_mie_q : _1740_;
  assign _1732_ = _1799_ ? \u_csr.u_csrfile.csr_mip_q : _1742_;
  assign _1735_ = _1799_ ? \u_csr.u_csrfile.csr_mtvec_q : _1745_;
  assign _1723_ = _1800_ ? 2'h0 : \u_csr.u_csrfile.csr_sr_q [12:11];
  assign _1744_ = _1799_ ? \u_csr.u_csrfile.csr_mtval_q : _1752_;
  assign _1762_ = _1799_ ? \u_csr.u_csrfile.csr_mcause_q : _1766_;
  assign _1739_ = _1799_ ? \u_csr.u_csrfile.csr_mepc_q : _1750_;
  assign \u_csr.u_csrfile.csr_sr_r [31:13] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [31:13] : _1769_[31:13];
  assign \u_csr.u_csrfile.csr_sr_r [10:9] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [10:9] : _1769_[10:9];
  assign \u_csr.u_csrfile.csr_sr_r [6] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [6] : _1769_[6];
  assign \u_csr.u_csrfile.csr_sr_r [4] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [4] : _1769_[4];
  assign \u_csr.u_csrfile.csr_sr_r [2] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [2] : _1769_[2];
  assign \u_csr.u_csrfile.csr_sr_r [0] = _1796_ ? \u_csr.u_csrfile.csr_sr_q [0] : _1769_[0];
  assign _1754_ = \u_csr.interrupt_w [11] ? 32'h8000000b : \u_csr.u_csrfile.csr_mcause_q ;
  assign _1749_ = \u_csr.interrupt_w [7] ? 32'h80000007 : _1754_;
  assign _1738_ = \u_csr.interrupt_w [3] ? 32'h80000003 : _1749_;
  assign _1729_ = _1797_ ? _1738_ : \u_csr.u_csrfile.csr_mcause_q ;
  assign _1734_ = _1797_ ? 32'h00000000 : \u_csr.u_csrfile.csr_mtval_q ;
  assign _1730_ = _1797_ ? \u_csr.u_csrfile.exception_pc_i : \u_csr.u_csrfile.csr_mepc_q ;
  assign _1746_ = _1797_ ? 1'h0 : \u_csr.u_csrfile.csr_sr_q [3];
  assign _1765_ = _1797_ ? \u_csr.u_csrfile.csr_mpriv_q : \u_csr.u_csrfile.csr_sr_q [12:11];
  assign _1759_[0] = _1797_ ? \u_csr.u_csrfile.csr_sr_q [3] : \u_csr.u_csrfile.csr_sr_q [7];
  assign _1759_[1] = _1797_ ? \u_csr.u_csrfile.csr_sr_q [8] : _1798_;
  assign _1753_ = _1797_ ? \u_csr.u_csrfile.csr_sr_q [5] : \u_csr.u_csrfile.csr_sr_q [1];
  assign _1736_ = _1797_ ? \u_csr.u_csrfile.csr_sr_q [1] : 1'h0;
  assign \u_csr.u_csrfile.csr_sr_r [12:11] = _1796_ ? _1765_ : _1769_[12:11];
  assign \u_csr.u_csrfile.csr_sr_r [8:7] = _1796_ ? _1759_ : _1769_[8:7];
  assign \u_csr.u_csrfile.csr_sr_r [5] = _1796_ ? _1753_ : _1769_[5];
  assign \u_csr.u_csrfile.csr_sr_r [3] = _1796_ ? _1746_ : _1769_[3];
  assign \u_csr.u_csrfile.csr_sr_r [1] = _1796_ ? _1736_ : _1769_[1];
  assign \u_csr.u_csrfile.csr_mtval_r = _1796_ ? _1734_ : _1744_;
  assign \u_csr.u_csrfile.csr_mcause_r = _1796_ ? _1729_ : _1762_;
  assign \u_csr.u_csrfile.csr_mepc_r = _1796_ ? _1730_ : _1739_;
  assign \u_csr.u_csrfile.csr_mscratch_r = _1796_ ? \u_csr.u_csrfile.csr_mscratch_q : _1733_;
  assign \u_csr.u_csrfile.csr_mie_r = _1796_ ? \u_csr.u_csrfile.csr_mie_q : _1731_;
  assign _1726_ = _1796_ ? \u_csr.u_csrfile.csr_mip_q : _1732_;
  assign \u_csr.u_csrfile.csr_mtvec_r = _1796_ ? \u_csr.u_csrfile.csr_mtvec_q : _1735_;
  logic [351:0] fangyuan22;
  assign fangyuan22 = { _1775_, _1776_, _1777_, _1778_, _1779_, _1780_, _1781_, _1782_, \u_csr.u_csrfile.csr_mcycle_q , cpu_id_i, 16'h4000, 16'h1100 };
  logic [10:0] fangyuan23;
  assign fangyuan23 = { _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1792_, _1837_, _1836_, _1834_, _1833_ };
  always @(32'h00000000 or fangyuan22 or fangyuan23) begin
    casez (fangyuan23)
      11'b??????????1 :
        \u_csr.csr_rdata_w = fangyuan22 [31:0] ;
      11'b?????????1? :
        \u_csr.csr_rdata_w = fangyuan22 [63:32] ;
      11'b????????1?? :
        \u_csr.csr_rdata_w = fangyuan22 [95:64] ;
      11'b???????1??? :
        \u_csr.csr_rdata_w = fangyuan22 [127:96] ;
      11'b??????1???? :
        \u_csr.csr_rdata_w = fangyuan22 [159:128] ;
      11'b?????1????? :
        \u_csr.csr_rdata_w = fangyuan22 [191:160] ;
      11'b????1?????? :
        \u_csr.csr_rdata_w = fangyuan22 [223:192] ;
      11'b???1??????? :
        \u_csr.csr_rdata_w = fangyuan22 [255:224] ;
      11'b??1???????? :
        \u_csr.csr_rdata_w = fangyuan22 [287:256] ;
      11'b?1????????? :
        \u_csr.csr_rdata_w = fangyuan22 [319:288] ;
      11'b1?????????? :
        \u_csr.csr_rdata_w = fangyuan22 [351:320] ;
      default:
        \u_csr.csr_rdata_w = 32'h00000000 ;
    endcase
  end
  assign _1833_ = \u_csr.opcode_opcode_i [31:20] == 10'h301;
  assign _1834_ = \u_csr.opcode_opcode_i [31:20] == 12'hf14;
  logic [1:0] fangyuan24;
  assign fangyuan24 = { _1835_[0], _1835_[1] };
  assign _1836_ = | fangyuan24;
  assign _1835_[0] = \u_csr.opcode_opcode_i [31:20] == 12'hc00;
  assign _1835_[1] = \u_csr.opcode_opcode_i [31:20] == 12'hc01;
  assign _1837_ = \u_csr.opcode_opcode_i [31:20] == 10'h304;
  assign _1838_ = \u_csr.opcode_opcode_i [31:20] == 10'h300;
  assign _1839_ = \u_csr.opcode_opcode_i [31:20] == 10'h343;
  assign _1840_ = \u_csr.opcode_opcode_i [31:20] == 10'h342;
  assign _1841_ = \u_csr.opcode_opcode_i [31:20] == 10'h305;
  assign _1842_ = \u_csr.opcode_opcode_i [31:20] == 10'h341;
  assign _1843_ = \u_csr.opcode_opcode_i [31:20] == 10'h340;
  assign _1844_ = _1813_ ? 1'h0 : \u_csr.u_csrfile.csr_mip_upd_q ;
  assign _1845_ = _1811_ ? 1'h1 : _1844_;
  assign _1715_ = rst_i ? 1'h0 : _1845_;
  assign _1846_ = _1847_ ? 2'h3 : \u_csr.u_csrfile.irq_priv_q ;
  assign _1720_ = rst_i ? 2'h3 : _1846_;
  logic [31:0] fangyuan25;
  assign fangyuan25 = { \u_csr.interrupt_w [0], \u_csr.interrupt_w [1], \u_csr.interrupt_w [2], \u_csr.interrupt_w [3], \u_csr.interrupt_w [4], \u_csr.interrupt_w [5], \u_csr.interrupt_w [6], \u_csr.interrupt_w [7], \u_csr.interrupt_w [8], \u_csr.interrupt_w [9], \u_csr.interrupt_w [10], \u_csr.interrupt_w [11], \u_csr.interrupt_w [12], \u_csr.interrupt_w [13], \u_csr.interrupt_w [14], \u_csr.interrupt_w [15], \u_csr.interrupt_w [16], \u_csr.interrupt_w [17], \u_csr.interrupt_w [18], \u_csr.interrupt_w [19], \u_csr.interrupt_w [20], \u_csr.interrupt_w [21], \u_csr.interrupt_w [22], \u_csr.interrupt_w [23], \u_csr.interrupt_w [24], \u_csr.interrupt_w [25], \u_csr.interrupt_w [26], \u_csr.interrupt_w [27], \u_csr.interrupt_w [28], \u_csr.interrupt_w [29], \u_csr.interrupt_w [30], \u_csr.interrupt_w [31] };
  assign _1847_ = | fangyuan25;
  logic [5:0] fangyuan26;
  assign fangyuan26 = { \u_csr.u_csrfile.exception_i [0], \u_csr.u_csrfile.exception_i [1], \u_csr.u_csrfile.exception_i [2], \u_csr.u_csrfile.exception_i [3], \u_csr.u_csrfile.exception_i [4], \u_csr.u_csrfile.exception_i [5] };
  assign _1848_ = | fangyuan26;
  assign \u_csr.interrupt_w = \u_csr.u_csrfile.csr_sr_q [3] ? \u_csr.u_csrfile.irq_pending_r : 32'h00000000;
  logic [31:0] fangyuan27;
  assign fangyuan27 = { \u_csr.u_csrfile.csr_mip_next_q [31:12], \u_csr.u_csrfile.csr_mip_next_r [11], \u_csr.u_csrfile.csr_mip_next_q [10], \u_csr.u_csrfile.csr_mip_next_r [9], \u_csr.u_csrfile.csr_mip_next_q [8], \u_csr.u_csrfile.csr_mip_next_r [7], \u_csr.u_csrfile.csr_mip_next_q [6], \u_csr.u_csrfile.csr_mip_next_r [5], \u_csr.u_csrfile.csr_mip_next_q [4:0] };
  assign _1849_ = \u_csr.u_csrfile.buffer_mip_w ? fangyuan27 : 32'h00000000;
  assign _1850_ = _1797_ ? \u_csr.u_csrfile.csr_mtvec_q : \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign _1866_ = \u_csr.opcode_opcode_i & 32'hfe00707f;
  assign \u_div.div_start_w = \u_div.opcode_valid_i & \u_div.div_rem_inst_w ;
  assign \u_div.div_complete_w = _1884_ & \u_div.div_busy_q ;
  assign _1867_ = \u_div.last_a_q == \u_csr.opcode_ra_operand_i ;
  assign _1868_ = \u_div.last_b_q == \u_div.opcode_rb_operand_i ;
  assign _1869_ = \u_div.last_div_q == \u_div.inst_div_w ;
  assign _1870_ = \u_div.last_divu_q == \u_div.inst_divu_w ;
  assign _1871_ = \u_div.last_rem_q == \u_div.inst_rem_w ;
  assign _1872_ = \u_div.last_remu_q == \u_div.inst_remu_w ;
  assign \u_div.inst_div_w = _1866_ == 26'h2004033;
  assign \u_div.inst_rem_w = _1866_ == 26'h2006033;
  assign \u_div.inst_divu_w = _1866_ == 26'h2005033;
  assign \u_div.inst_remu_w = _1866_ == 26'h2007033;
  assign _1873_ = \u_div.divisor_q <= \u_div.dividend_q ;
  assign _1874_ = _1867_ && _1868_;
  assign _1875_ = _1874_ && _1869_;
  assign _1876_ = _1875_ && _1870_;
  assign _1877_ = _1876_ && _1871_;
  assign _1878_ = _1877_ && _1872_;
  assign _1879_ = \u_div.signed_operation_w && \u_csr.opcode_ra_operand_i [31];
  assign _1880_ = \u_div.signed_operation_w && \u_div.opcode_rb_operand_i [31];
  assign _1881_ = \u_div.inst_div_w && _1887_;
  assign _1882_ = _1881_ && _1932_;
  assign _1883_ = \u_div.inst_rem_w && \u_csr.opcode_ra_operand_i [31];
  assign _1884_ = ! _1933_;
  assign _1885_ = _1882_ || _1883_;
  assign \u_div.div_operation_w = \u_div.inst_div_w || \u_div.inst_divu_w ;
  assign _1886_ = \u_div.div_operation_w || \u_div.inst_rem_w ;
  assign \u_div.div_rem_inst_w = _1886_ || \u_div.inst_remu_w ;
  assign \u_div.signed_operation_w = \u_div.inst_div_w || \u_div.inst_rem_w ;
  assign _1887_ = \u_csr.opcode_ra_operand_i [31] != \u_div.opcode_rb_operand_i [31];
  assign _1888_ = - \u_csr.opcode_ra_operand_i ;
  assign _1889_ = - \u_div.opcode_rb_operand_i ;
  assign _1890_ = - \u_div.quotient_q ;
  assign _1891_ = - \u_div.dividend_q ;
  assign _1892_ = \u_div.quotient_q | \u_div.q_mask_q ;
  always @(posedge clk_i)
      \u_div.wb_result_q <= _1865_;
  always @(posedge clk_i)
      \u_div.valid_q <= _1864_;
  always @(posedge clk_i)
      \u_div.dividend_q <= _1853_;
  always @(posedge clk_i)
      \u_div.divisor_q <= _1854_;
  always @(posedge clk_i)
      \u_div.quotient_q <= _1863_;
  always @(posedge clk_i)
      \u_div.q_mask_q <= _1862_;
  always @(posedge clk_i)
      \u_div.div_inst_q <= _1852_;
  always @(posedge clk_i)
      \u_div.div_busy_q <= _1851_;
  always @(posedge clk_i)
      \u_div.invert_res_q <= _1855_;
  always @(posedge clk_i)
      \u_div.last_a_q <= _1856_;
  always @(posedge clk_i)
      \u_div.last_b_q <= _1857_;
  always @(posedge clk_i)
      \u_div.last_div_q <= _1858_;
  always @(posedge clk_i)
      \u_div.last_divu_q <= _1859_;
  always @(posedge clk_i)
      \u_div.last_rem_q <= _1860_;
  always @(posedge clk_i)
      \u_div.last_remu_q <= _1861_;
  assign _1893_ = \u_div.div_complete_w ? \u_div.div_result_r : \u_div.wb_result_q ;
  assign _1865_ = rst_i ? 32'h00000000 : _1893_;
  assign _1864_ = rst_i ? 1'h0 : \u_div.div_complete_w ;
  assign \u_div.div_result_r = \u_div.div_inst_q ? _1935_ : _1936_;
  assign _1894_ = _1878_ ? \u_div.last_remu_q : \u_div.inst_remu_w ;
  assign _1895_ = \u_div.div_start_w ? _1894_ : \u_div.last_remu_q ;
  assign _1861_ = rst_i ? 1'h0 : _1895_;
  assign _1896_ = _1878_ ? \u_div.last_rem_q : \u_div.inst_rem_w ;
  assign _1897_ = \u_div.div_start_w ? _1896_ : \u_div.last_rem_q ;
  assign _1860_ = rst_i ? 1'h0 : _1897_;
  assign _1898_ = _1878_ ? \u_div.last_divu_q : \u_div.inst_divu_w ;
  assign _1899_ = \u_div.div_start_w ? _1898_ : \u_div.last_divu_q ;
  assign _1859_ = rst_i ? 1'h0 : _1899_;
  assign _1900_ = _1878_ ? \u_div.last_div_q : \u_div.inst_div_w ;
  assign _1901_ = \u_div.div_start_w ? _1900_ : \u_div.last_div_q ;
  assign _1858_ = rst_i ? 1'h0 : _1901_;
  assign _1902_ = _1878_ ? \u_div.last_b_q : \u_div.opcode_rb_operand_i ;
  assign _1903_ = \u_div.div_start_w ? _1902_ : \u_div.last_b_q ;
  assign _1857_ = rst_i ? 32'h00000000 : _1903_;
  assign _1904_ = _1878_ ? \u_div.last_a_q : \u_csr.opcode_ra_operand_i ;
  assign _1905_ = \u_div.div_start_w ? _1904_ : \u_div.last_a_q ;
  assign _1856_ = rst_i ? 32'h00000000 : _1905_;
  assign _1906_ = _1878_ ? \u_div.invert_res_q : _1885_;
  assign _1907_ = \u_div.div_start_w ? _1906_ : \u_div.invert_res_q ;
  assign _1855_ = rst_i ? 1'h0 : _1907_;
  assign _1908_ = \u_div.div_complete_w ? 1'h0 : \u_div.div_busy_q ;
  assign _1909_ = \u_div.div_start_w ? 1'h1 : _1908_;
  assign _1851_ = rst_i ? 1'h0 : _1909_;
  assign _1910_ = _1878_ ? \u_div.div_inst_q : \u_div.div_operation_w ;
  assign _1911_ = \u_div.div_start_w ? _1910_ : \u_div.div_inst_q ;
  assign _1852_ = rst_i ? 1'h0 : _1911_;
  logic [31:0] fangyuan28;
  assign fangyuan28 = { 1'h0, \u_div.q_mask_q [31:1] };
  assign _1912_ = \u_div.div_busy_q ? fangyuan28 : \u_div.q_mask_q ;
  assign _1913_ = \u_div.div_complete_w ? \u_div.q_mask_q : _1912_;
  assign _1914_ = _1878_ ? \u_div.q_mask_q : 32'h80000000;
  assign _1915_ = \u_div.div_start_w ? _1914_ : _1913_;
  assign _1862_ = rst_i ? 32'h00000000 : _1915_;
  assign _1916_ = _1873_ ? _1892_ : \u_div.quotient_q ;
  assign _1917_ = \u_div.div_busy_q ? _1916_ : \u_div.quotient_q ;
  assign _1918_ = \u_div.div_complete_w ? \u_div.quotient_q : _1917_;
  assign _1919_ = _1878_ ? \u_div.quotient_q : 32'h00000000;
  assign _1920_ = \u_div.div_start_w ? _1919_ : _1918_;
  assign _1863_ = rst_i ? 32'h00000000 : _1920_;
  logic [62:0] fangyuan29;
  assign fangyuan29 = { 1'h0, \u_div.divisor_q [62:1] };
  assign _1921_ = \u_div.div_busy_q ? fangyuan29 : \u_div.divisor_q ;
  assign _1922_ = \u_div.div_complete_w ? \u_div.divisor_q : _1921_;
  logic [62:0] fangyuan30;
  assign fangyuan30 = { _1889_, 16'h0000, 15'h0000 };
  logic [62:0] fangyuan31;
  assign fangyuan31 = { \u_div.opcode_rb_operand_i , 16'h0000, 15'h0000 };
  assign _1923_ = _1880_ ? fangyuan30 : fangyuan31;
  assign _1924_ = _1878_ ? \u_div.divisor_q : _1923_;
  assign _1925_ = \u_div.div_start_w ? _1924_ : _1922_;
  assign _1854_ = rst_i ? 63'h0000000000000000 : _1925_;
  assign _1926_ = _1873_ ? _1934_ : \u_div.dividend_q ;
  assign _1927_ = \u_div.div_busy_q ? _1926_ : \u_div.dividend_q ;
  assign _1928_ = \u_div.div_complete_w ? \u_div.dividend_q : _1927_;
  assign _1929_ = _1879_ ? _1888_ : \u_csr.opcode_ra_operand_i ;
  assign _1930_ = _1878_ ? \u_div.dividend_q : _1929_;
  assign _1931_ = \u_div.div_start_w ? _1930_ : _1928_;
  assign _1853_ = rst_i ? 32'h00000000 : _1931_;
  logic [31:0] fangyuan32;
  assign fangyuan32 = { \u_div.opcode_rb_operand_i [0], \u_div.opcode_rb_operand_i [1], \u_div.opcode_rb_operand_i [2], \u_div.opcode_rb_operand_i [3], \u_div.opcode_rb_operand_i [4], \u_div.opcode_rb_operand_i [5], \u_div.opcode_rb_operand_i [6], \u_div.opcode_rb_operand_i [7], \u_div.opcode_rb_operand_i [8], \u_div.opcode_rb_operand_i [9], \u_div.opcode_rb_operand_i [10], \u_div.opcode_rb_operand_i [11], \u_div.opcode_rb_operand_i [12], \u_div.opcode_rb_operand_i [13], \u_div.opcode_rb_operand_i [14], \u_div.opcode_rb_operand_i [15], \u_div.opcode_rb_operand_i [16], \u_div.opcode_rb_operand_i [17], \u_div.opcode_rb_operand_i [18], \u_div.opcode_rb_operand_i [19], \u_div.opcode_rb_operand_i [20], \u_div.opcode_rb_operand_i [21], \u_div.opcode_rb_operand_i [22], \u_div.opcode_rb_operand_i [23], \u_div.opcode_rb_operand_i [24], \u_div.opcode_rb_operand_i [25], \u_div.opcode_rb_operand_i [26], \u_div.opcode_rb_operand_i [27], \u_div.opcode_rb_operand_i [28], \u_div.opcode_rb_operand_i [29], \u_div.opcode_rb_operand_i [30], \u_div.opcode_rb_operand_i [31] };
  assign _1932_ = | fangyuan32;
  logic [31:0] fangyuan33;
  assign fangyuan33 = { \u_div.q_mask_q [0], \u_div.q_mask_q [1], \u_div.q_mask_q [2], \u_div.q_mask_q [3], \u_div.q_mask_q [4], \u_div.q_mask_q [5], \u_div.q_mask_q [6], \u_div.q_mask_q [7], \u_div.q_mask_q [8], \u_div.q_mask_q [9], \u_div.q_mask_q [10], \u_div.q_mask_q [11], \u_div.q_mask_q [12], \u_div.q_mask_q [13], \u_div.q_mask_q [14], \u_div.q_mask_q [15], \u_div.q_mask_q [16], \u_div.q_mask_q [17], \u_div.q_mask_q [18], \u_div.q_mask_q [19], \u_div.q_mask_q [20], \u_div.q_mask_q [21], \u_div.q_mask_q [22], \u_div.q_mask_q [23], \u_div.q_mask_q [24], \u_div.q_mask_q [25], \u_div.q_mask_q [26], \u_div.q_mask_q [27], \u_div.q_mask_q [28], \u_div.q_mask_q [29], \u_div.q_mask_q [30], \u_div.q_mask_q [31] };
  assign _1933_ = | fangyuan33;
  assign _1934_ = \u_div.dividend_q - \u_div.divisor_q [31:0];
  assign _1935_ = \u_div.invert_res_q ? _1890_ : \u_div.quotient_q ;
  assign _1936_ = \u_div.invert_res_q ? _1891_ : \u_div.dividend_q ;
  logic [31:0] fangyuan34;
  assign fangyuan34 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [7], \u_csr.opcode_opcode_i [30:25], \u_csr.opcode_opcode_i [11:8], 1'h0 };
  assign _2027_ = \u_exec0.opcode_pc_i + fangyuan34;
  logic [31:0] fangyuan35;
  assign fangyuan35 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [19:12], \u_csr.opcode_opcode_i [20], \u_csr.opcode_opcode_i [30:21], 1'h0 };
  assign _2028_ = \u_exec0.opcode_pc_i + fangyuan35;
  logic [31:0] fangyuan36;
  assign fangyuan36 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _2029_ = \u_csr.opcode_ra_operand_i + fangyuan36;
  assign _2030_ = \u_exec0.opcode_pc_i + 3'h4;
  assign _2031_ = \u_csr.opcode_opcode_i & 32'hfe00707f;
  assign _2032_ = \u_csr.opcode_opcode_i & 15'h707f;
  assign _2033_ = \u_csr.opcode_opcode_i & 32'hfc00707f;
  assign _2034_ = \u_csr.opcode_opcode_i & 7'h7f;
  assign _2035_ = \u_div.opcode_valid_i & \u_exec0.branch_taken_r ;
  assign _2036_ = \u_div.opcode_valid_i & _2085_;
  assign _2037_ = _2031_ == 15'h7033;
  assign _2038_ = _2031_ == 15'h6033;
  assign _2039_ = _2031_ == 13'h1033;
  assign _2040_ = _2031_ == 31'h40005033;
  assign _2041_ = _2031_ == 15'h5033;
  assign _2042_ = _2031_ == 31'h40000033;
  assign _2043_ = _2031_ == 15'h4033;
  assign _2044_ = _2031_ == 14'h2033;
  assign _2045_ = _2031_ == 14'h3033;
  assign _2046_ = _2032_ == 5'h13;
  assign _2047_ = _2032_ == 15'h7013;
  assign _2048_ = _2032_ == 14'h2013;
  assign _2049_ = _2032_ == 14'h3013;
  assign _2050_ = _2032_ == 15'h6013;
  assign _2051_ = _2032_ == 15'h4013;
  assign _2052_ = _2033_ == 13'h1013;
  assign _2053_ = _2033_ == 15'h5013;
  assign _2054_ = _2033_ == 31'h40005013;
  assign _2055_ = _2034_ == 6'h37;
  assign _2056_ = _2034_ == 5'h17;
  assign _2057_ = _2034_ == 7'h6f;
  assign _2058_ = _2032_ == 7'h67;
  assign _2059_ = \u_csr.opcode_opcode_i [11:7] == 1'h1;
  assign _2060_ = \u_csr.opcode_opcode_i [19:15] == 1'h1;
  assign _2061_ = ! \u_csr.opcode_opcode_i [31:20];
  assign _2062_ = _2032_ == 7'h63;
  assign _2063_ = \u_csr.opcode_ra_operand_i == \u_div.opcode_rb_operand_i ;
  assign _2064_ = _2032_ == 13'h1063;
  assign _2065_ = _2032_ == 15'h4063;
  assign _2066_ = _2032_ == 15'h5063;
  assign _2067_ = _2032_ == 15'h6063;
  assign _2068_ = _2032_ == 15'h7063;
  assign _2069_ = _2031_ == 6'h33;
  assign _2070_ = \u_csr.opcode_ra_operand_i >= \u_div.opcode_rb_operand_i ;
  assign _2071_ = _2060_ && _2061_;
  assign _2072_ = _2083_ && _2059_;
  assign _2073_ = \u_exec0.branch_r && _2035_;
  assign _2074_ = \u_exec0.branch_r && _2036_;
  assign _2075_ = \u_exec0.branch_r && \u_div.opcode_valid_i ;
  assign _2076_ = _2075_ && \u_exec0.branch_call_r ;
  assign _2077_ = _2075_ && \u_exec0.branch_ret_r ;
  assign _2078_ = _2075_ && \u_exec0.branch_jmp_r ;
  assign \u_exec0.branch_d_request_o = _2075_ && \u_exec0.branch_taken_r ;
  assign _2079_ = _2057_ || _2058_;
  assign _2080_ = \u_csr.opcode_ra_operand_i < \u_div.opcode_rb_operand_i ;
  assign _2081_ = \u_csr.opcode_ra_operand_i [31] != \u_div.opcode_rb_operand_i [31];
  assign _2082_ = \u_csr.opcode_ra_operand_i != \u_div.opcode_rb_operand_i ;
  assign _2083_ = ~ _2071_;
  assign _2084_ = ~ _2086_;
  assign _2085_ = ~ \u_exec0.branch_taken_r ;
  assign _2086_ = _2072_ | _2071_;
  assign _2087_ = _2013_ | _2063_;
  always @(posedge clk_i)
      \u_exec0.branch_taken_q <= _1941_;
  always @(posedge clk_i)
      \u_exec0.branch_ntaken_q <= _1939_;
  always @(posedge clk_i)
      \u_exec0.pc_x_q <= _1943_;
  always @(posedge clk_i)
      \u_exec0.pc_m_q <= _1942_;
  always @(posedge clk_i)
      \u_exec0.branch_call_q <= _1937_;
  always @(posedge clk_i)
      \u_exec0.branch_ret_q <= _1940_;
  always @(posedge clk_i)
      \u_exec0.branch_jmp_q <= _1938_;
  always @(posedge clk_i)
      \u_exec0.result_q <= _1944_;
  assign _2088_ = \u_div.opcode_valid_i ? _2078_ : \u_exec0.branch_jmp_q ;
  assign _1938_ = rst_i ? 1'h0 : _2088_;
  assign _2089_ = \u_div.opcode_valid_i ? _2077_ : \u_exec0.branch_ret_q ;
  assign _1940_ = rst_i ? 1'h0 : _2089_;
  assign _2090_ = \u_div.opcode_valid_i ? _2076_ : \u_exec0.branch_call_q ;
  assign _1937_ = rst_i ? 1'h0 : _2090_;
  assign _2091_ = \u_div.opcode_valid_i ? \u_exec0.opcode_pc_i : \u_exec0.pc_m_q ;
  assign _1942_ = rst_i ? 32'h00000000 : _2091_;
  assign _2092_ = \u_div.opcode_valid_i ? _2098_ : \u_exec0.pc_x_q ;
  assign _1943_ = rst_i ? 32'h00000000 : _2092_;
  assign _2093_ = \u_div.opcode_valid_i ? _2074_ : \u_exec0.branch_ntaken_q ;
  assign _1939_ = rst_i ? 1'h0 : _2093_;
  assign _2094_ = \u_div.opcode_valid_i ? _2073_ : \u_exec0.branch_taken_q ;
  assign _1941_ = rst_i ? 1'h0 : _2094_;
  assign _2023_ = _2068_ ? _2070_ : 1'h0;
  assign _2022_ = _2068_ ? 1'h1 : 1'h0;
  assign _2018_ = _2067_ ? _2080_ : _2023_;
  assign _2017_ = _2067_ ? 1'h1 : _2022_;
  assign _2013_ = _2081_ ? \u_div.opcode_rb_operand_i [31] : _2097_[31];
  assign _2012_ = _2066_ ? _2087_ : _2018_;
  assign _2011_ = _2066_ ? 1'h1 : _2017_;
  assign _2007_ = _2081_ ? \u_csr.opcode_ra_operand_i [31] : _2096_[31];
  assign _2006_ = _2065_ ? _2007_ : _2012_;
  assign _2005_ = _2065_ ? 1'h1 : _2011_;
  assign _2001_ = _2064_ ? _2082_ : _2006_;
  assign _2000_ = _2064_ ? 1'h1 : _2005_;
  assign _1996_ = _2062_ ? _2063_ : _2001_;
  assign _1995_ = _2062_ ? 1'h1 : _2000_;
  assign _1991_[31:1] = _2058_ ? _2029_[31:1] : _2027_[31:1];
  assign _1986_ = _2058_ ? _2072_ : 1'h0;
  assign _1989_ = _2058_ ? _2071_ : 1'h0;
  assign _1987_ = _2058_ ? _2084_ : 1'h0;
  assign _1991_[0] = _2058_ ? 1'h0 : _2027_[0];
  assign _1990_ = _2058_ ? 1'h1 : _1996_;
  assign _1988_ = _2058_ ? 1'h1 : _1995_;
  assign \u_exec0.branch_jmp_r = _2057_ ? 1'h1 : _1987_;
  assign \u_exec0.branch_call_r = _2057_ ? _2059_ : _1986_;
  assign \u_exec0.branch_target_r = _2057_ ? _2028_ : _1991_;
  assign \u_exec0.branch_taken_r = _2057_ ? 1'h1 : _1990_;
  assign \u_exec0.branch_r = _2057_ ? 1'h1 : _1988_;
  assign \u_exec0.branch_ret_r = _2057_ ? 1'h0 : _1989_;
  assign _2095_ = \u_exec0.hold_i ? \u_exec0.result_q : \u_exec0.alu_p_w ;
  assign _1944_ = rst_i ? 32'h00000000 : _2095_;
  assign _1981_ = _2079_ ? 3'h4 : 3'h0;
  assign _1982_ = _2079_ ? \u_exec0.opcode_pc_i : 32'h00000000;
  logic [31:0] fangyuan37;
  assign fangyuan37 = { \u_csr.opcode_opcode_i [31:12], 12'h000 };
  logic [31:0] fangyuan38;
  assign fangyuan38 = { 29'h00000000, _1981_ };
  assign _1980_ = _2056_ ? fangyuan37 : fangyuan38;
  assign _1979_ = _2056_ ? \u_exec0.opcode_pc_i : _1982_;
  logic [3:0] fangyuan39;
  assign fangyuan39 = { 1'h0, _1981_ };
  assign _1978_ = _2056_ ? 4'h4 : fangyuan39;
  logic [31:0] fangyuan40;
  assign fangyuan40 = { \u_csr.opcode_opcode_i [31:12], 12'h000 };
  assign _1976_ = _2055_ ? fangyuan40 : _1979_;
  assign _1977_ = _2055_ ? 32'h00000000 : _1980_;
  assign _1975_ = _2055_ ? 4'h0 : _1978_;
  logic [31:0] fangyuan41;
  assign fangyuan41 = { 27'h0000000, \u_csr.opcode_opcode_i [24:20] };
  assign _1974_ = _2054_ ? fangyuan41 : _1977_;
  assign _1973_ = _2054_ ? \u_csr.opcode_ra_operand_i : _1976_;
  assign _1972_ = _2054_ ? 4'h3 : _1975_;
  logic [31:0] fangyuan42;
  assign fangyuan42 = { 27'h0000000, \u_csr.opcode_opcode_i [24:20] };
  assign _1971_ = _2053_ ? fangyuan42 : _1974_;
  assign _1970_ = _2053_ ? \u_csr.opcode_ra_operand_i : _1973_;
  assign _1969_ = _2053_ ? 4'h2 : _1972_;
  logic [31:0] fangyuan43;
  assign fangyuan43 = { 27'h0000000, \u_csr.opcode_opcode_i [24:20] };
  assign _1968_ = _2052_ ? fangyuan43 : _1971_;
  assign _1967_ = _2052_ ? \u_csr.opcode_ra_operand_i : _1970_;
  assign _1966_ = _2052_ ? 4'h1 : _1969_;
  logic [31:0] fangyuan44;
  assign fangyuan44 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1965_ = _2051_ ? fangyuan44 : _1968_;
  assign _1964_ = _2051_ ? \u_csr.opcode_ra_operand_i : _1967_;
  assign _1963_ = _2051_ ? 4'h9 : _1966_;
  logic [31:0] fangyuan45;
  assign fangyuan45 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1962_ = _2050_ ? fangyuan45 : _1965_;
  assign _1961_ = _2050_ ? \u_csr.opcode_ra_operand_i : _1964_;
  assign _1960_ = _2050_ ? 4'h8 : _1963_;
  logic [31:0] fangyuan46;
  assign fangyuan46 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1959_ = _2049_ ? fangyuan46 : _1962_;
  assign _1958_ = _2049_ ? \u_csr.opcode_ra_operand_i : _1961_;
  assign _1957_ = _2049_ ? 4'ha : _1960_;
  logic [31:0] fangyuan47;
  assign fangyuan47 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1956_ = _2048_ ? fangyuan47 : _1959_;
  assign _1955_ = _2048_ ? \u_csr.opcode_ra_operand_i : _1958_;
  assign _1954_ = _2048_ ? 4'hb : _1957_;
  logic [31:0] fangyuan48;
  assign fangyuan48 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1953_ = _2047_ ? fangyuan48 : _1956_;
  assign _1952_ = _2047_ ? \u_csr.opcode_ra_operand_i : _1955_;
  assign _1951_ = _2047_ ? 4'h7 : _1954_;
  logic [31:0] fangyuan49;
  assign fangyuan49 = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign _1950_ = _2046_ ? fangyuan49 : _1953_;
  assign _1949_ = _2046_ ? \u_csr.opcode_ra_operand_i : _1952_;
  assign _1948_ = _2046_ ? 4'h4 : _1951_;
  assign _1947_ = _2045_ ? \u_div.opcode_rb_operand_i : _1950_;
  assign _1946_ = _2045_ ? \u_csr.opcode_ra_operand_i : _1949_;
  assign _1945_ = _2045_ ? 4'ha : _1948_;
  assign _2026_ = _2044_ ? \u_div.opcode_rb_operand_i : _1947_;
  assign _2025_ = _2044_ ? \u_csr.opcode_ra_operand_i : _1946_;
  assign _2024_ = _2044_ ? 4'hb : _1945_;
  assign _2021_ = _2043_ ? \u_div.opcode_rb_operand_i : _2026_;
  assign _2020_ = _2043_ ? \u_csr.opcode_ra_operand_i : _2025_;
  assign _2019_ = _2043_ ? 4'h9 : _2024_;
  assign _2016_ = _2042_ ? \u_div.opcode_rb_operand_i : _2021_;
  assign _2015_ = _2042_ ? \u_csr.opcode_ra_operand_i : _2020_;
  assign _2014_ = _2042_ ? 4'h6 : _2019_;
  assign _2010_ = _2041_ ? \u_div.opcode_rb_operand_i : _2016_;
  assign _2009_ = _2041_ ? \u_csr.opcode_ra_operand_i : _2015_;
  assign _2008_ = _2041_ ? 4'h2 : _2014_;
  assign _2004_ = _2040_ ? \u_div.opcode_rb_operand_i : _2010_;
  assign _2003_ = _2040_ ? \u_csr.opcode_ra_operand_i : _2009_;
  assign _2002_ = _2040_ ? 4'h3 : _2008_;
  assign _1999_ = _2039_ ? \u_div.opcode_rb_operand_i : _2004_;
  assign _1998_ = _2039_ ? \u_csr.opcode_ra_operand_i : _2003_;
  assign _1997_ = _2039_ ? 4'h1 : _2002_;
  assign _1994_ = _2038_ ? \u_div.opcode_rb_operand_i : _1999_;
  assign _1993_ = _2038_ ? \u_csr.opcode_ra_operand_i : _1998_;
  assign _1992_ = _2038_ ? 4'h8 : _1997_;
  assign _1985_ = _2037_ ? \u_div.opcode_rb_operand_i : _1994_;
  assign _1984_ = _2037_ ? \u_csr.opcode_ra_operand_i : _1993_;
  assign _1983_ = _2037_ ? 4'h7 : _1992_;
  assign \u_exec0.alu_input_b_r = _2069_ ? \u_div.opcode_rb_operand_i : _1985_;
  assign \u_exec0.alu_input_a_r = _2069_ ? \u_csr.opcode_ra_operand_i : _1984_;
  assign \u_exec0.alu_func_r = _2069_ ? 4'h4 : _1983_;
  assign _2096_ = \u_csr.opcode_ra_operand_i - \u_div.opcode_rb_operand_i ;
  assign _2097_ = \u_div.opcode_rb_operand_i - \u_csr.opcode_ra_operand_i ;
  assign _2098_ = \u_exec0.branch_taken_r ? \u_exec0.branch_target_r : _2030_;
  assign _2111_ = \u_exec0.alu_input_a_r + \u_exec0.alu_input_b_r ;
  assign _2112_ = \u_exec0.alu_input_a_r & \u_exec0.alu_input_b_r ;
  assign _2115_ = \u_exec0.alu_func_r == 2'h3;
  assign _2116_ = \u_exec0.alu_input_a_r [31] && _2115_;
  assign _2117_ = \u_exec0.alu_input_a_r < \u_exec0.alu_input_b_r ;
  assign _2118_ = \u_exec0.alu_input_a_r [31] != \u_exec0.alu_input_b_r [31];
  assign _2119_ = \u_exec0.alu_input_a_r | \u_exec0.alu_input_b_r ;
  assign _2110_ = _2118_ ? _2129_[0] : _2130_[0];
  assign _2120_ = \u_exec0.alu_func_r == 4'hb;
  logic [31:0] fangyuan50;
  assign fangyuan50 = { _2108_, _2107_[31:16] };
  assign _2109_ = \u_exec0.alu_input_b_r [4] ? fangyuan50 : _2107_;
  assign _2113_[0] = \u_exec0.alu_func_r == 2'h2;
  logic [31:0] fangyuan51;
  assign fangyuan51 = { _2108_[15:8], _2106_[31:8] };
  assign _2107_ = \u_exec0.alu_input_b_r [3] ? fangyuan51 : _2106_;
  logic [31:0] fangyuan52;
  assign fangyuan52 = { _2108_[15:12], _2105_[31:4] };
  assign _2106_ = \u_exec0.alu_input_b_r [2] ? fangyuan52 : _2105_;
  logic [1:0] fangyuan53;
  assign fangyuan53 = { _2115_, _2113_[0] };
  assign _2121_ = | fangyuan53;
  logic [31:0] fangyuan54;
  assign fangyuan54 = { _2108_[15:14], _2104_[31:2] };
  assign _2105_ = \u_exec0.alu_input_b_r [1] ? fangyuan54 : _2104_;
  logic [31:0] fangyuan55;
  assign fangyuan55 = { _2108_[15], \u_exec0.alu_input_a_r [31:1] };
  assign _2104_ = \u_exec0.alu_input_b_r [0] ? fangyuan55 : \u_exec0.alu_input_a_r ;
  assign _2108_ = _2116_ ? 16'hffff : 16'h0000;
  logic [31:0] fangyuan56;
  assign fangyuan56 = { _2103_[15:0], 16'h0000 };
  assign _2099_ = \u_exec0.alu_input_b_r [4] ? fangyuan56 : _2103_;
  assign _2122_ = \u_exec0.alu_func_r == 1'h1;
  logic [31:0] fangyuan57;
  assign fangyuan57 = { _2102_[23:0], 8'h00 };
  assign _2103_ = \u_exec0.alu_input_b_r [3] ? fangyuan57 : _2102_;
  logic [31:0] fangyuan58;
  assign fangyuan58 = { _2101_[27:0], 4'h0 };
  assign _2102_ = \u_exec0.alu_input_b_r [2] ? fangyuan58 : _2101_;
  logic [31:0] fangyuan59;
  assign fangyuan59 = { _2100_[29:0], 2'h0 };
  assign _2101_ = \u_exec0.alu_input_b_r [1] ? fangyuan59 : _2100_;
  logic [31:0] fangyuan60;
  assign fangyuan60 = { \u_exec0.alu_input_a_r [30:0], 1'h0 };
  assign _2100_ = \u_exec0.alu_input_b_r [0] ? fangyuan60 : \u_exec0.alu_input_a_r ;
  logic [287:0] fangyuan61;
  assign fangyuan61 = { _2099_, _2109_, _2111_, \u_exec0.u_alu.sub_res_w , _2112_, _2119_, _2131_, 16'h0000, 15'h0000, _2114_[0], 16'h0000, 15'h0000, _2110_ };
  logic [8:0] fangyuan62;
  assign fangyuan62 = { _2122_, _2121_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2120_ };
  always @(\u_exec0.alu_input_a_r or fangyuan61 or fangyuan62) begin
    casez (fangyuan62)
      9'b????????1 :
        \u_exec0.alu_p_w = fangyuan61 [31:0] ;
      9'b???????1? :
        \u_exec0.alu_p_w = fangyuan61 [63:32] ;
      9'b??????1?? :
        \u_exec0.alu_p_w = fangyuan61 [95:64] ;
      9'b?????1??? :
        \u_exec0.alu_p_w = fangyuan61 [127:96] ;
      9'b????1???? :
        \u_exec0.alu_p_w = fangyuan61 [159:128] ;
      9'b???1????? :
        \u_exec0.alu_p_w = fangyuan61 [191:160] ;
      9'b??1?????? :
        \u_exec0.alu_p_w = fangyuan61 [223:192] ;
      9'b?1??????? :
        \u_exec0.alu_p_w = fangyuan61 [255:224] ;
      9'b1???????? :
        \u_exec0.alu_p_w = fangyuan61 [287:256] ;
      default:
        \u_exec0.alu_p_w = \u_exec0.alu_input_a_r ;
    endcase
  end
  assign _2123_ = \u_exec0.alu_func_r == 4'ha;
  assign _2124_ = \u_exec0.alu_func_r == 4'h9;
  assign _2125_ = \u_exec0.alu_func_r == 4'h8;
  assign _2126_ = \u_exec0.alu_func_r == 3'h7;
  assign _2127_ = \u_exec0.alu_func_r == 3'h6;
  assign _2128_ = \u_exec0.alu_func_r == 3'h4;
  assign \u_exec0.u_alu.sub_res_w = \u_exec0.alu_input_a_r - \u_exec0.alu_input_b_r ;
  assign _2114_[0] = _2117_ ? 1'h1 : 1'h0;
  assign _2129_[0] = \u_exec0.alu_input_a_r [31] ? 1'h1 : 1'h0;
  assign _2130_[0] = \u_exec0.u_alu.sub_res_w [31] ? 1'h1 : 1'h0;
  assign _2131_ = \u_exec0.alu_input_a_r ^ \u_exec0.alu_input_b_r ;
  logic [31:0] fangyuan63;
  assign fangyuan63 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [7], \u_exec1.opcode_opcode_i [30:25], \u_exec1.opcode_opcode_i [11:8], 1'h0 };
  assign _2222_ = \u_exec1.opcode_pc_i + fangyuan63;
  logic [31:0] fangyuan64;
  assign fangyuan64 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [19:12], \u_exec1.opcode_opcode_i [20], \u_exec1.opcode_opcode_i [30:21], 1'h0 };
  assign _2223_ = \u_exec1.opcode_pc_i + fangyuan64;
  logic [31:0] fangyuan65;
  assign fangyuan65 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2224_ = \u_exec1.opcode_ra_operand_i + fangyuan65;
  assign _2225_ = \u_exec1.opcode_pc_i + 3'h4;
  assign _2226_ = \u_exec1.opcode_opcode_i & 32'hfe00707f;
  assign _2227_ = \u_exec1.opcode_opcode_i & 15'h707f;
  assign _2228_ = \u_exec1.opcode_opcode_i & 32'hfc00707f;
  assign _2229_ = \u_exec1.opcode_opcode_i & 7'h7f;
  assign _2230_ = \u_exec1.opcode_valid_i & \u_exec1.branch_taken_r ;
  assign _2231_ = \u_exec1.opcode_valid_i & _2280_;
  assign _2232_ = _2226_ == 15'h7033;
  assign _2233_ = _2226_ == 15'h6033;
  assign _2234_ = _2226_ == 13'h1033;
  assign _2235_ = _2226_ == 31'h40005033;
  assign _2236_ = _2226_ == 15'h5033;
  assign _2237_ = _2226_ == 31'h40000033;
  assign _2238_ = _2226_ == 15'h4033;
  assign _2239_ = _2226_ == 14'h2033;
  assign _2240_ = _2226_ == 14'h3033;
  assign _2241_ = _2227_ == 5'h13;
  assign _2242_ = _2227_ == 15'h7013;
  assign _2243_ = _2227_ == 14'h2013;
  assign _2244_ = _2227_ == 14'h3013;
  assign _2245_ = _2227_ == 15'h6013;
  assign _2246_ = _2227_ == 15'h4013;
  assign _2247_ = _2228_ == 13'h1013;
  assign _2248_ = _2228_ == 15'h5013;
  assign _2249_ = _2228_ == 31'h40005013;
  assign _2250_ = _2229_ == 6'h37;
  assign _2251_ = _2229_ == 5'h17;
  assign _2252_ = _2229_ == 7'h6f;
  assign _2253_ = _2227_ == 7'h67;
  assign _2254_ = \u_exec1.opcode_opcode_i [11:7] == 1'h1;
  assign _2255_ = \u_exec1.opcode_opcode_i [19:15] == 1'h1;
  assign _2256_ = ! \u_exec1.opcode_opcode_i [31:20];
  assign _2257_ = _2227_ == 7'h63;
  assign _2258_ = \u_exec1.opcode_ra_operand_i == \u_exec1.opcode_rb_operand_i ;
  assign _2259_ = _2227_ == 13'h1063;
  assign _2260_ = _2227_ == 15'h4063;
  assign _2261_ = _2227_ == 15'h5063;
  assign _2262_ = _2227_ == 15'h6063;
  assign _2263_ = _2227_ == 15'h7063;
  assign _2264_ = _2226_ == 6'h33;
  assign _2265_ = \u_exec1.opcode_ra_operand_i >= \u_exec1.opcode_rb_operand_i ;
  assign _2266_ = _2255_ && _2256_;
  assign _2267_ = _2278_ && _2254_;
  assign _2268_ = \u_exec1.branch_r && _2230_;
  assign _2269_ = \u_exec1.branch_r && _2231_;
  assign _2270_ = \u_exec1.branch_r && \u_exec1.opcode_valid_i ;
  assign _2271_ = _2270_ && \u_exec1.branch_call_r ;
  assign _2272_ = _2270_ && \u_exec1.branch_ret_r ;
  assign _2273_ = _2270_ && \u_exec1.branch_jmp_r ;
  assign \u_exec1.branch_d_request_o = _2270_ && \u_exec1.branch_taken_r ;
  assign _2274_ = _2252_ || _2253_;
  assign _2275_ = \u_exec1.opcode_ra_operand_i < \u_exec1.opcode_rb_operand_i ;
  assign _2276_ = \u_exec1.opcode_ra_operand_i [31] != \u_exec1.opcode_rb_operand_i [31];
  assign _2277_ = \u_exec1.opcode_ra_operand_i != \u_exec1.opcode_rb_operand_i ;
  assign _2278_ = ~ _2266_;
  assign _2279_ = ~ _2281_;
  assign _2280_ = ~ \u_exec1.branch_taken_r ;
  assign _2281_ = _2267_ | _2266_;
  assign _2282_ = _2208_ | _2258_;
  assign \u_exec1.branch_request_o = \u_exec1.branch_taken_q | \u_exec1.branch_ntaken_q ;
  always @(posedge clk_i)
      \u_exec1.branch_taken_q <= _2136_;
  always @(posedge clk_i)
      \u_exec1.branch_ntaken_q <= _2134_;
  always @(posedge clk_i)
      \u_exec1.pc_x_q <= _2138_;
  always @(posedge clk_i)
      \u_exec1.pc_m_q <= _2137_;
  always @(posedge clk_i)
      \u_exec1.branch_call_q <= _2132_;
  always @(posedge clk_i)
      \u_exec1.branch_ret_q <= _2135_;
  always @(posedge clk_i)
      \u_exec1.branch_jmp_q <= _2133_;
  always @(posedge clk_i)
      \u_exec1.result_q <= _2139_;
  assign _2283_ = \u_exec1.opcode_valid_i ? _2273_ : \u_exec1.branch_jmp_q ;
  assign _2133_ = rst_i ? 1'h0 : _2283_;
  assign _2284_ = \u_exec1.opcode_valid_i ? _2272_ : \u_exec1.branch_ret_q ;
  assign _2135_ = rst_i ? 1'h0 : _2284_;
  assign _2285_ = \u_exec1.opcode_valid_i ? _2271_ : \u_exec1.branch_call_q ;
  assign _2132_ = rst_i ? 1'h0 : _2285_;
  assign _2286_ = \u_exec1.opcode_valid_i ? \u_exec1.opcode_pc_i : \u_exec1.pc_m_q ;
  assign _2137_ = rst_i ? 32'h00000000 : _2286_;
  assign _2287_ = \u_exec1.opcode_valid_i ? _2293_ : \u_exec1.pc_x_q ;
  assign _2138_ = rst_i ? 32'h00000000 : _2287_;
  assign _2288_ = \u_exec1.opcode_valid_i ? _2269_ : \u_exec1.branch_ntaken_q ;
  assign _2134_ = rst_i ? 1'h0 : _2288_;
  assign _2289_ = \u_exec1.opcode_valid_i ? _2268_ : \u_exec1.branch_taken_q ;
  assign _2136_ = rst_i ? 1'h0 : _2289_;
  assign _2218_ = _2263_ ? _2265_ : 1'h0;
  assign _2217_ = _2263_ ? 1'h1 : 1'h0;
  assign _2213_ = _2262_ ? _2275_ : _2218_;
  assign _2212_ = _2262_ ? 1'h1 : _2217_;
  assign _2208_ = _2276_ ? \u_exec1.opcode_rb_operand_i [31] : _2292_[31];
  assign _2207_ = _2261_ ? _2282_ : _2213_;
  assign _2206_ = _2261_ ? 1'h1 : _2212_;
  assign _2202_ = _2276_ ? \u_exec1.opcode_ra_operand_i [31] : _2291_[31];
  assign _2201_ = _2260_ ? _2202_ : _2207_;
  assign _2200_ = _2260_ ? 1'h1 : _2206_;
  assign _2196_ = _2259_ ? _2277_ : _2201_;
  assign _2195_ = _2259_ ? 1'h1 : _2200_;
  assign _2191_ = _2257_ ? _2258_ : _2196_;
  assign _2190_ = _2257_ ? 1'h1 : _2195_;
  assign _2186_[31:1] = _2253_ ? _2224_[31:1] : _2222_[31:1];
  assign _2181_ = _2253_ ? _2267_ : 1'h0;
  assign _2184_ = _2253_ ? _2266_ : 1'h0;
  assign _2182_ = _2253_ ? _2279_ : 1'h0;
  assign _2186_[0] = _2253_ ? 1'h0 : _2222_[0];
  assign _2185_ = _2253_ ? 1'h1 : _2191_;
  assign _2183_ = _2253_ ? 1'h1 : _2190_;
  assign \u_exec1.branch_jmp_r = _2252_ ? 1'h1 : _2182_;
  assign \u_exec1.branch_call_r = _2252_ ? _2254_ : _2181_;
  assign \u_exec1.branch_target_r = _2252_ ? _2223_ : _2186_;
  assign \u_exec1.branch_taken_r = _2252_ ? 1'h1 : _2185_;
  assign \u_exec1.branch_r = _2252_ ? 1'h1 : _2183_;
  assign \u_exec1.branch_ret_r = _2252_ ? 1'h0 : _2184_;
  assign _2290_ = \u_exec0.hold_i ? \u_exec1.result_q : \u_exec1.alu_p_w ;
  assign _2139_ = rst_i ? 32'h00000000 : _2290_;
  assign _2176_ = _2274_ ? 3'h4 : 3'h0;
  assign _2177_ = _2274_ ? \u_exec1.opcode_pc_i : 32'h00000000;
  logic [31:0] fangyuan66;
  assign fangyuan66 = { \u_exec1.opcode_opcode_i [31:12], 12'h000 };
  logic [31:0] fangyuan67;
  assign fangyuan67 = { 29'h00000000, _2176_ };
  assign _2175_ = _2251_ ? fangyuan66 : fangyuan67;
  assign _2174_ = _2251_ ? \u_exec1.opcode_pc_i : _2177_;
  logic [3:0] fangyuan68;
  assign fangyuan68 = { 1'h0, _2176_ };
  assign _2173_ = _2251_ ? 4'h4 : fangyuan68;
  logic [31:0] fangyuan69;
  assign fangyuan69 = { \u_exec1.opcode_opcode_i [31:12], 12'h000 };
  assign _2171_ = _2250_ ? fangyuan69 : _2174_;
  assign _2172_ = _2250_ ? 32'h00000000 : _2175_;
  assign _2170_ = _2250_ ? 4'h0 : _2173_;
  logic [31:0] fangyuan70;
  assign fangyuan70 = { 27'h0000000, \u_exec1.opcode_opcode_i [24:20] };
  assign _2169_ = _2249_ ? fangyuan70 : _2172_;
  assign _2168_ = _2249_ ? \u_exec1.opcode_ra_operand_i : _2171_;
  assign _2167_ = _2249_ ? 4'h3 : _2170_;
  logic [31:0] fangyuan71;
  assign fangyuan71 = { 27'h0000000, \u_exec1.opcode_opcode_i [24:20] };
  assign _2166_ = _2248_ ? fangyuan71 : _2169_;
  assign _2165_ = _2248_ ? \u_exec1.opcode_ra_operand_i : _2168_;
  assign _2164_ = _2248_ ? 4'h2 : _2167_;
  logic [31:0] fangyuan72;
  assign fangyuan72 = { 27'h0000000, \u_exec1.opcode_opcode_i [24:20] };
  assign _2163_ = _2247_ ? fangyuan72 : _2166_;
  assign _2162_ = _2247_ ? \u_exec1.opcode_ra_operand_i : _2165_;
  assign _2161_ = _2247_ ? 4'h1 : _2164_;
  logic [31:0] fangyuan73;
  assign fangyuan73 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2160_ = _2246_ ? fangyuan73 : _2163_;
  assign _2159_ = _2246_ ? \u_exec1.opcode_ra_operand_i : _2162_;
  assign _2158_ = _2246_ ? 4'h9 : _2161_;
  logic [31:0] fangyuan74;
  assign fangyuan74 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2157_ = _2245_ ? fangyuan74 : _2160_;
  assign _2156_ = _2245_ ? \u_exec1.opcode_ra_operand_i : _2159_;
  assign _2155_ = _2245_ ? 4'h8 : _2158_;
  logic [31:0] fangyuan75;
  assign fangyuan75 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2154_ = _2244_ ? fangyuan75 : _2157_;
  assign _2153_ = _2244_ ? \u_exec1.opcode_ra_operand_i : _2156_;
  assign _2152_ = _2244_ ? 4'ha : _2155_;
  logic [31:0] fangyuan76;
  assign fangyuan76 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2151_ = _2243_ ? fangyuan76 : _2154_;
  assign _2150_ = _2243_ ? \u_exec1.opcode_ra_operand_i : _2153_;
  assign _2149_ = _2243_ ? 4'hb : _2152_;
  logic [31:0] fangyuan77;
  assign fangyuan77 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2148_ = _2242_ ? fangyuan77 : _2151_;
  assign _2147_ = _2242_ ? \u_exec1.opcode_ra_operand_i : _2150_;
  assign _2146_ = _2242_ ? 4'h7 : _2149_;
  logic [31:0] fangyuan78;
  assign fangyuan78 = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign _2145_ = _2241_ ? fangyuan78 : _2148_;
  assign _2144_ = _2241_ ? \u_exec1.opcode_ra_operand_i : _2147_;
  assign _2143_ = _2241_ ? 4'h4 : _2146_;
  assign _2142_ = _2240_ ? \u_exec1.opcode_rb_operand_i : _2145_;
  assign _2141_ = _2240_ ? \u_exec1.opcode_ra_operand_i : _2144_;
  assign _2140_ = _2240_ ? 4'ha : _2143_;
  assign _2221_ = _2239_ ? \u_exec1.opcode_rb_operand_i : _2142_;
  assign _2220_ = _2239_ ? \u_exec1.opcode_ra_operand_i : _2141_;
  assign _2219_ = _2239_ ? 4'hb : _2140_;
  assign _2216_ = _2238_ ? \u_exec1.opcode_rb_operand_i : _2221_;
  assign _2215_ = _2238_ ? \u_exec1.opcode_ra_operand_i : _2220_;
  assign _2214_ = _2238_ ? 4'h9 : _2219_;
  assign _2211_ = _2237_ ? \u_exec1.opcode_rb_operand_i : _2216_;
  assign _2210_ = _2237_ ? \u_exec1.opcode_ra_operand_i : _2215_;
  assign _2209_ = _2237_ ? 4'h6 : _2214_;
  assign _2205_ = _2236_ ? \u_exec1.opcode_rb_operand_i : _2211_;
  assign _2204_ = _2236_ ? \u_exec1.opcode_ra_operand_i : _2210_;
  assign _2203_ = _2236_ ? 4'h2 : _2209_;
  assign _2199_ = _2235_ ? \u_exec1.opcode_rb_operand_i : _2205_;
  assign _2198_ = _2235_ ? \u_exec1.opcode_ra_operand_i : _2204_;
  assign _2197_ = _2235_ ? 4'h3 : _2203_;
  assign _2194_ = _2234_ ? \u_exec1.opcode_rb_operand_i : _2199_;
  assign _2193_ = _2234_ ? \u_exec1.opcode_ra_operand_i : _2198_;
  assign _2192_ = _2234_ ? 4'h1 : _2197_;
  assign _2189_ = _2233_ ? \u_exec1.opcode_rb_operand_i : _2194_;
  assign _2188_ = _2233_ ? \u_exec1.opcode_ra_operand_i : _2193_;
  assign _2187_ = _2233_ ? 4'h8 : _2192_;
  assign _2180_ = _2232_ ? \u_exec1.opcode_rb_operand_i : _2189_;
  assign _2179_ = _2232_ ? \u_exec1.opcode_ra_operand_i : _2188_;
  assign _2178_ = _2232_ ? 4'h7 : _2187_;
  assign \u_exec1.alu_input_b_r = _2264_ ? \u_exec1.opcode_rb_operand_i : _2180_;
  assign \u_exec1.alu_input_a_r = _2264_ ? \u_exec1.opcode_ra_operand_i : _2179_;
  assign \u_exec1.alu_func_r = _2264_ ? 4'h4 : _2178_;
  assign _2291_ = \u_exec1.opcode_ra_operand_i - \u_exec1.opcode_rb_operand_i ;
  assign _2292_ = \u_exec1.opcode_rb_operand_i - \u_exec1.opcode_ra_operand_i ;
  assign _2293_ = \u_exec1.branch_taken_r ? \u_exec1.branch_target_r : _2225_;
  assign _2306_ = \u_exec1.alu_input_a_r + \u_exec1.alu_input_b_r ;
  assign _2307_ = \u_exec1.alu_input_a_r & \u_exec1.alu_input_b_r ;
  assign _2310_ = \u_exec1.alu_func_r == 2'h3;
  assign _2311_ = \u_exec1.alu_input_a_r [31] && _2310_;
  assign _2312_ = \u_exec1.alu_input_a_r < \u_exec1.alu_input_b_r ;
  assign _2313_ = \u_exec1.alu_input_a_r [31] != \u_exec1.alu_input_b_r [31];
  assign _2314_ = \u_exec1.alu_input_a_r | \u_exec1.alu_input_b_r ;
  assign _2305_ = _2313_ ? _2324_[0] : _2325_[0];
  assign _2315_ = \u_exec1.alu_func_r == 4'hb;
  logic [31:0] fangyuan79;
  assign fangyuan79 = { _2303_, _2302_[31:16] };
  assign _2304_ = \u_exec1.alu_input_b_r [4] ? fangyuan79 : _2302_;
  assign _2308_[0] = \u_exec1.alu_func_r == 2'h2;
  logic [31:0] fangyuan80;
  assign fangyuan80 = { _2303_[15:8], _2301_[31:8] };
  assign _2302_ = \u_exec1.alu_input_b_r [3] ? fangyuan80 : _2301_;
  logic [31:0] fangyuan81;
  assign fangyuan81 = { _2303_[15:12], _2300_[31:4] };
  assign _2301_ = \u_exec1.alu_input_b_r [2] ? fangyuan81 : _2300_;
  logic [1:0] fangyuan82;
  assign fangyuan82 = { _2310_, _2308_[0] };
  assign _2316_ = | fangyuan82;
  logic [31:0] fangyuan83;
  assign fangyuan83 = { _2303_[15:14], _2299_[31:2] };
  assign _2300_ = \u_exec1.alu_input_b_r [1] ? fangyuan83 : _2299_;
  logic [31:0] fangyuan84;
  assign fangyuan84 = { _2303_[15], \u_exec1.alu_input_a_r [31:1] };
  assign _2299_ = \u_exec1.alu_input_b_r [0] ? fangyuan84 : \u_exec1.alu_input_a_r ;
  assign _2303_ = _2311_ ? 16'hffff : 16'h0000;
  logic [31:0] fangyuan85;
  assign fangyuan85 = { _2298_[15:0], 16'h0000 };
  assign _2294_ = \u_exec1.alu_input_b_r [4] ? fangyuan85 : _2298_;
  assign _2317_ = \u_exec1.alu_func_r == 1'h1;
  logic [31:0] fangyuan86;
  assign fangyuan86 = { _2297_[23:0], 8'h00 };
  assign _2298_ = \u_exec1.alu_input_b_r [3] ? fangyuan86 : _2297_;
  logic [31:0] fangyuan87;
  assign fangyuan87 = { _2296_[27:0], 4'h0 };
  assign _2297_ = \u_exec1.alu_input_b_r [2] ? fangyuan87 : _2296_;
  logic [31:0] fangyuan88;
  assign fangyuan88 = { _2295_[29:0], 2'h0 };
  assign _2296_ = \u_exec1.alu_input_b_r [1] ? fangyuan88 : _2295_;
  logic [31:0] fangyuan89;
  assign fangyuan89 = { \u_exec1.alu_input_a_r [30:0], 1'h0 };
  assign _2295_ = \u_exec1.alu_input_b_r [0] ? fangyuan89 : \u_exec1.alu_input_a_r ;
  logic [287:0] fangyuan90;
  assign fangyuan90 = { _2294_, _2304_, _2306_, \u_exec1.u_alu.sub_res_w , _2307_, _2314_, _2326_, 16'h0000, 15'h0000, _2309_[0], 16'h0000, 15'h0000, _2305_ };
  logic [8:0] fangyuan91;
  assign fangyuan91 = { _2317_, _2316_, _2323_, _2322_, _2321_, _2320_, _2319_, _2318_, _2315_ };
  always @(\u_exec1.alu_input_a_r or fangyuan90 or fangyuan91) begin
    casez (fangyuan91)
      9'b????????1 :
        \u_exec1.alu_p_w = fangyuan90 [31:0] ;
      9'b???????1? :
        \u_exec1.alu_p_w = fangyuan90 [63:32] ;
      9'b??????1?? :
        \u_exec1.alu_p_w = fangyuan90 [95:64] ;
      9'b?????1??? :
        \u_exec1.alu_p_w = fangyuan90 [127:96] ;
      9'b????1???? :
        \u_exec1.alu_p_w = fangyuan90 [159:128] ;
      9'b???1????? :
        \u_exec1.alu_p_w = fangyuan90 [191:160] ;
      9'b??1?????? :
        \u_exec1.alu_p_w = fangyuan90 [223:192] ;
      9'b?1??????? :
        \u_exec1.alu_p_w = fangyuan90 [255:224] ;
      9'b1???????? :
        \u_exec1.alu_p_w = fangyuan90 [287:256] ;
      default:
        \u_exec1.alu_p_w = \u_exec1.alu_input_a_r ;
    endcase
  end
  assign _2318_ = \u_exec1.alu_func_r == 4'ha;
  assign _2319_ = \u_exec1.alu_func_r == 4'h9;
  assign _2320_ = \u_exec1.alu_func_r == 4'h8;
  assign _2321_ = \u_exec1.alu_func_r == 3'h7;
  assign _2322_ = \u_exec1.alu_func_r == 3'h6;
  assign _2323_ = \u_exec1.alu_func_r == 3'h4;
  assign \u_exec1.u_alu.sub_res_w = \u_exec1.alu_input_a_r - \u_exec1.alu_input_b_r ;
  assign _2309_[0] = _2312_ ? 1'h1 : 1'h0;
  assign _2324_[0] = \u_exec1.alu_input_a_r [31] ? 1'h1 : 1'h0;
  assign _2325_[0] = \u_exec1.u_alu.sub_res_w [31] ? 1'h1 : 1'h0;
  assign _2326_ = \u_exec1.alu_input_a_r ^ \u_exec1.alu_input_b_r ;
  assign _2327_ = \u_frontend.u_decode.fetch_in_fault_page_i | \u_frontend.u_decode.fetch_in_fault_fetch_i ;
  assign \u_frontend.u_decode.u_dec0.fetch_fault_i = \u_frontend.u_decode.u_fifo.info0_out_o [0] | \u_frontend.u_decode.u_fifo.info0_out_o [1];
  assign \u_frontend.u_decode.u_dec1.fetch_fault_i = \u_frontend.u_decode.u_fifo.info1_out_o [0] | \u_frontend.u_decode.u_fifo.info1_out_o [1];
  assign \u_frontend.u_decode.u_fifo.data_in_i = _2327_ ? 64'h0000000000000000 : \u_frontend.u_decode.fetch_in_instr_i ;
  assign _2328_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hfe00707f;
  assign _2329_ = \u_frontend.u_decode.u_fifo.data0_out_o & 15'h707f;
  assign _2330_ = \u_frontend.u_decode.u_fifo.data0_out_o & 7'h7f;
  assign _2331_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hfc00707f;
  assign _2332_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hffffffff;
  assign _2333_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hdfffffff;
  assign _2334_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hffff8fff;
  assign _2335_ = \u_frontend.u_decode.u_fifo.data0_out_o & 32'hfe007fff;
  assign _2336_ = _2328_ == 26'h2003033;
  assign _2337_ = _2328_ == 26'h2004033;
  assign _2338_ = _2328_ == 26'h2005033;
  assign _2339_ = _2328_ == 26'h2006033;
  assign _2340_ = _2328_ == 26'h2007033;
  assign _2341_ = _2329_ == 7'h67;
  assign _2342_ = _2330_ == 7'h6f;
  assign _2343_ = _2330_ == 6'h37;
  assign _2344_ = _2330_ == 5'h17;
  assign _2345_ = _2329_ == 5'h13;
  assign _2346_ = _2331_ == 13'h1013;
  assign _2347_ = _2329_ == 14'h2013;
  assign _2348_ = _2329_ == 14'h3013;
  assign _2349_ = _2329_ == 15'h4013;
  assign _2350_ = _2331_ == 15'h5013;
  assign _2351_ = _2331_ == 31'h40005013;
  assign _2352_ = _2329_ == 15'h6013;
  assign _2353_ = _2329_ == 15'h7013;
  assign _2354_ = _2328_ == 6'h33;
  assign _2355_ = _2328_ == 31'h40000033;
  assign _2356_ = _2328_ == 13'h1033;
  assign _2357_ = _2328_ == 14'h2033;
  assign _2358_ = _2328_ == 14'h3033;
  assign _2359_ = _2328_ == 15'h4033;
  assign _2360_ = _2328_ == 15'h5033;
  assign _2361_ = _2328_ == 31'h40005033;
  assign _2362_ = _2328_ == 15'h6033;
  assign _2363_ = _2328_ == 15'h7033;
  assign _2364_ = _2329_ == 2'h3;
  assign _2365_ = _2329_ == 13'h1003;
  assign _2366_ = _2329_ == 14'h2003;
  assign _2367_ = _2329_ == 15'h4003;
  assign _2368_ = _2329_ == 15'h5003;
  assign _2369_ = _2329_ == 15'h6003;
  assign _2370_ = _2328_ == 26'h2000033;
  assign _2371_ = _2328_ == 26'h2001033;
  assign _2372_ = _2328_ == 26'h2002033;
  assign _2373_ = _2329_ == 13'h1073;
  assign _2374_ = _2329_ == 14'h2073;
  assign _2375_ = _2329_ == 14'h3073;
  assign _2376_ = _2329_ == 15'h5073;
  assign _2377_ = _2329_ == 15'h6073;
  assign _2378_ = _2329_ == 15'h7073;
  assign _2379_ = _2329_ == 6'h23;
  assign _2380_ = _2329_ == 13'h1023;
  assign _2381_ = _2329_ == 14'h2023;
  assign _2382_ = _2329_ == 7'h63;
  assign _2383_ = _2329_ == 13'h1063;
  assign _2384_ = _2329_ == 15'h4063;
  assign _2385_ = _2329_ == 15'h5063;
  assign _2386_ = _2329_ == 15'h6063;
  assign _2387_ = _2329_ == 15'h7063;
  assign _2388_ = _2332_ == 7'h73;
  assign _2389_ = _2332_ == 21'h100073;
  assign _2390_ = _2333_ == 29'h10200073;
  assign _2391_ = _2334_ == 29'h10500073;
  assign _2392_ = _2329_ == 4'hf;
  assign _2393_ = _2329_ == 13'h100f;
  assign _2394_ = _2335_ == 29'h12000073;
  assign _2395_ = 1'h1 && _2336_;
  assign _2396_ = 1'h1 && _2337_;
  assign _2397_ = 1'h1 && _2338_;
  assign _2398_ = 1'h1 && _2339_;
  assign _2399_ = 1'h1 && _2340_;
  assign \u_frontend.u_decode.u_dec0.invalid_w = \u_frontend.u_decode.u_dec0.valid_i && _2532_;
  assign \u_frontend.u_decode.u_dec0.mul_o = 1'h1 && _2482_;
  assign \u_frontend.u_decode.u_dec0.div_o = 1'h1 && _2485_;
  assign _2400_ = 1'h1 && _2370_;
  assign _2401_ = 1'h1 && _2371_;
  assign _2402_ = 1'h1 && _2372_;
  assign _2403_ = _2531_ || _2395_;
  assign _2404_ = _2403_ || _2396_;
  assign _2405_ = _2404_ || _2397_;
  assign _2406_ = _2405_ || _2398_;
  assign _2407_ = _2406_ || _2399_;
  assign _2408_ = _2341_ || _2342_;
  assign _2409_ = _2408_ || _2343_;
  assign _2410_ = _2409_ || _2344_;
  assign _2411_ = _2410_ || _2345_;
  assign _2412_ = _2411_ || _2346_;
  assign _2413_ = _2412_ || _2347_;
  assign _2414_ = _2413_ || _2348_;
  assign _2415_ = _2414_ || _2349_;
  assign _2416_ = _2415_ || _2350_;
  assign _2417_ = _2416_ || _2351_;
  assign _2418_ = _2417_ || _2352_;
  assign _2419_ = _2418_ || _2353_;
  assign _2420_ = _2419_ || _2354_;
  assign _2421_ = _2420_ || _2355_;
  assign _2422_ = _2421_ || _2356_;
  assign _2423_ = _2422_ || _2357_;
  assign _2424_ = _2423_ || _2358_;
  assign _2425_ = _2424_ || _2359_;
  assign _2426_ = _2425_ || _2360_;
  assign _2427_ = _2426_ || _2361_;
  assign _2428_ = _2427_ || _2362_;
  assign _2429_ = _2428_ || _2363_;
  assign _2430_ = _2429_ || _2364_;
  assign _2431_ = _2430_ || _2365_;
  assign _2432_ = _2431_ || _2366_;
  assign _2433_ = _2432_ || _2367_;
  assign _2434_ = _2433_ || _2368_;
  assign _2435_ = _2434_ || _2369_;
  assign _2436_ = _2435_ || _2370_;
  assign _2437_ = _2436_ || _2371_;
  assign _2438_ = _2437_ || _2372_;
  assign _2439_ = _2438_ || _2336_;
  assign _2440_ = _2439_ || _2337_;
  assign _2441_ = _2440_ || _2338_;
  assign _2442_ = _2441_ || _2339_;
  assign _2443_ = _2442_ || _2340_;
  assign _2444_ = _2443_ || _2373_;
  assign _2445_ = _2444_ || _2374_;
  assign _2446_ = _2445_ || _2375_;
  assign _2447_ = _2446_ || _2376_;
  assign _2448_ = _2447_ || _2377_;
  assign \u_frontend.u_decode.u_dec0.rd_valid_o = _2448_ || _2378_;
  assign _2449_ = _2353_ || _2345_;
  assign _2450_ = _2449_ || _2347_;
  assign _2451_ = _2450_ || _2348_;
  assign _2452_ = _2451_ || _2352_;
  assign _2453_ = _2452_ || _2349_;
  assign _2454_ = _2453_ || _2346_;
  assign _2455_ = _2454_ || _2350_;
  assign _2456_ = _2455_ || _2351_;
  assign _2457_ = _2456_ || _2343_;
  assign _2458_ = _2457_ || _2344_;
  assign _2459_ = _2458_ || _2354_;
  assign _2460_ = _2459_ || _2355_;
  assign _2461_ = _2460_ || _2357_;
  assign _2462_ = _2461_ || _2358_;
  assign _2463_ = _2462_ || _2359_;
  assign _2464_ = _2463_ || _2362_;
  assign _2465_ = _2464_ || _2363_;
  assign _2466_ = _2465_ || _2356_;
  assign _2467_ = _2466_ || _2360_;
  assign \u_frontend.u_decode.u_dec0.exec_o = _2467_ || _2361_;
  assign _2468_ = _2364_ || _2365_;
  assign _2469_ = _2468_ || _2366_;
  assign _2470_ = _2469_ || _2367_;
  assign _2471_ = _2470_ || _2368_;
  assign _2472_ = _2471_ || _2369_;
  assign _2473_ = _2472_ || _2379_;
  assign _2474_ = _2473_ || _2380_;
  assign \u_frontend.u_decode.u_dec0.lsu_o = _2474_ || _2381_;
  assign _2475_ = _2408_ || _2382_;
  assign _2476_ = _2475_ || _2383_;
  assign _2477_ = _2476_ || _2384_;
  assign _2478_ = _2477_ || _2385_;
  assign _2479_ = _2478_ || _2386_;
  assign \u_frontend.u_decode.u_dec0.branch_o = _2479_ || _2387_;
  assign _2480_ = _2370_ || _2371_;
  assign _2481_ = _2480_ || _2372_;
  assign _2482_ = _2481_ || _2336_;
  assign _2483_ = _2337_ || _2338_;
  assign _2484_ = _2483_ || _2339_;
  assign _2485_ = _2484_ || _2340_;
  assign _2486_ = _2388_ || _2389_;
  assign _2487_ = _2486_ || _2390_;
  assign _2488_ = _2487_ || _2373_;
  assign _2489_ = _2488_ || _2374_;
  assign _2490_ = _2489_ || _2375_;
  assign _2491_ = _2490_ || _2376_;
  assign _2492_ = _2491_ || _2377_;
  assign _2493_ = _2492_ || _2378_;
  assign _2494_ = _2493_ || _2391_;
  assign _2495_ = _2494_ || _2392_;
  assign _2496_ = _2495_ || _2393_;
  assign _2497_ = _2496_ || _2394_;
  assign _2498_ = _2497_ || \u_frontend.u_decode.u_dec0.invalid_w ;
  assign \u_frontend.u_decode.u_dec0.csr_o = _2498_ || \u_frontend.u_decode.u_dec0.fetch_fault_i ;
  assign _2499_ = \u_frontend.u_decode.u_dec0.exec_o || _2342_;
  assign _2500_ = _2499_ || _2341_;
  assign _2501_ = _2500_ || _2382_;
  assign _2502_ = _2501_ || _2383_;
  assign _2503_ = _2502_ || _2384_;
  assign _2504_ = _2503_ || _2385_;
  assign _2505_ = _2504_ || _2386_;
  assign _2506_ = _2505_ || _2387_;
  assign _2507_ = _2506_ || _2364_;
  assign _2508_ = _2507_ || _2365_;
  assign _2509_ = _2508_ || _2366_;
  assign _2510_ = _2509_ || _2367_;
  assign _2511_ = _2510_ || _2368_;
  assign _2512_ = _2511_ || _2369_;
  assign _2513_ = _2512_ || _2379_;
  assign _2514_ = _2513_ || _2380_;
  assign _2515_ = _2514_ || _2381_;
  assign _2516_ = _2515_ || _2388_;
  assign _2517_ = _2516_ || _2389_;
  assign _2518_ = _2517_ || _2390_;
  assign _2519_ = _2518_ || _2373_;
  assign _2520_ = _2519_ || _2374_;
  assign _2521_ = _2520_ || _2375_;
  assign _2522_ = _2521_ || _2376_;
  assign _2523_ = _2522_ || _2377_;
  assign _2524_ = _2523_ || _2378_;
  assign _2525_ = _2524_ || _2391_;
  assign _2526_ = _2525_ || _2392_;
  assign _2527_ = _2526_ || _2393_;
  assign _2528_ = _2527_ || _2394_;
  assign _2529_ = _2528_ || _2400_;
  assign _2530_ = _2529_ || _2401_;
  assign _2531_ = _2530_ || _2402_;
  assign _2532_ = ~ _2407_;
  assign _2533_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hfe00707f;
  assign _2534_ = \u_frontend.u_decode.u_fifo.data1_out_o & 15'h707f;
  assign _2535_ = \u_frontend.u_decode.u_fifo.data1_out_o & 7'h7f;
  assign _2536_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hfc00707f;
  assign _2537_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hffffffff;
  assign _2538_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hdfffffff;
  assign _2539_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hffff8fff;
  assign _2540_ = \u_frontend.u_decode.u_fifo.data1_out_o & 32'hfe007fff;
  assign _2541_ = _2533_ == 26'h2003033;
  assign _2542_ = _2533_ == 26'h2004033;
  assign _2543_ = _2533_ == 26'h2005033;
  assign _2544_ = _2533_ == 26'h2006033;
  assign _2545_ = _2533_ == 26'h2007033;
  assign _2546_ = _2534_ == 7'h67;
  assign _2547_ = _2535_ == 7'h6f;
  assign _2548_ = _2535_ == 6'h37;
  assign _2549_ = _2535_ == 5'h17;
  assign _2550_ = _2534_ == 5'h13;
  assign _2551_ = _2536_ == 13'h1013;
  assign _2552_ = _2534_ == 14'h2013;
  assign _2553_ = _2534_ == 14'h3013;
  assign _2554_ = _2534_ == 15'h4013;
  assign _2555_ = _2536_ == 15'h5013;
  assign _2556_ = _2536_ == 31'h40005013;
  assign _2557_ = _2534_ == 15'h6013;
  assign _2558_ = _2534_ == 15'h7013;
  assign _2559_ = _2533_ == 6'h33;
  assign _2560_ = _2533_ == 31'h40000033;
  assign _2561_ = _2533_ == 13'h1033;
  assign _2562_ = _2533_ == 14'h2033;
  assign _2563_ = _2533_ == 14'h3033;
  assign _2564_ = _2533_ == 15'h4033;
  assign _2565_ = _2533_ == 15'h5033;
  assign _2566_ = _2533_ == 31'h40005033;
  assign _2567_ = _2533_ == 15'h6033;
  assign _2568_ = _2533_ == 15'h7033;
  assign _2569_ = _2534_ == 2'h3;
  assign _2570_ = _2534_ == 13'h1003;
  assign _2571_ = _2534_ == 14'h2003;
  assign _2572_ = _2534_ == 15'h4003;
  assign _2573_ = _2534_ == 15'h5003;
  assign _2574_ = _2534_ == 15'h6003;
  assign _2575_ = _2533_ == 26'h2000033;
  assign _2576_ = _2533_ == 26'h2001033;
  assign _2577_ = _2533_ == 26'h2002033;
  assign _2578_ = _2534_ == 13'h1073;
  assign _2579_ = _2534_ == 14'h2073;
  assign _2580_ = _2534_ == 14'h3073;
  assign _2581_ = _2534_ == 15'h5073;
  assign _2582_ = _2534_ == 15'h6073;
  assign _2583_ = _2534_ == 15'h7073;
  assign _2584_ = _2534_ == 6'h23;
  assign _2585_ = _2534_ == 13'h1023;
  assign _2586_ = _2534_ == 14'h2023;
  assign _2587_ = _2534_ == 7'h63;
  assign _2588_ = _2534_ == 13'h1063;
  assign _2589_ = _2534_ == 15'h4063;
  assign _2590_ = _2534_ == 15'h5063;
  assign _2591_ = _2534_ == 15'h6063;
  assign _2592_ = _2534_ == 15'h7063;
  assign _2593_ = _2537_ == 7'h73;
  assign _2594_ = _2537_ == 21'h100073;
  assign _2595_ = _2538_ == 29'h10200073;
  assign _2596_ = _2539_ == 29'h10500073;
  assign _2597_ = _2534_ == 4'hf;
  assign _2598_ = _2534_ == 13'h100f;
  assign _2599_ = _2540_ == 29'h12000073;
  assign _2600_ = 1'h1 && _2541_;
  assign _2601_ = 1'h1 && _2542_;
  assign _2602_ = 1'h1 && _2543_;
  assign _2603_ = 1'h1 && _2544_;
  assign _2604_ = 1'h1 && _2545_;
  assign \u_frontend.u_decode.u_dec1.invalid_w = \u_frontend.u_decode.u_dec1.valid_i && _2737_;
  assign \u_frontend.u_decode.u_dec1.mul_o = 1'h1 && _2687_;
  assign \u_frontend.u_decode.u_dec1.div_o = 1'h1 && _2690_;
  assign _2605_ = 1'h1 && _2575_;
  assign _2606_ = 1'h1 && _2576_;
  assign _2607_ = 1'h1 && _2577_;
  assign _2608_ = _2736_ || _2600_;
  assign _2609_ = _2608_ || _2601_;
  assign _2610_ = _2609_ || _2602_;
  assign _2611_ = _2610_ || _2603_;
  assign _2612_ = _2611_ || _2604_;
  assign _2613_ = _2546_ || _2547_;
  assign _2614_ = _2613_ || _2548_;
  assign _2615_ = _2614_ || _2549_;
  assign _2616_ = _2615_ || _2550_;
  assign _2617_ = _2616_ || _2551_;
  assign _2618_ = _2617_ || _2552_;
  assign _2619_ = _2618_ || _2553_;
  assign _2620_ = _2619_ || _2554_;
  assign _2621_ = _2620_ || _2555_;
  assign _2622_ = _2621_ || _2556_;
  assign _2623_ = _2622_ || _2557_;
  assign _2624_ = _2623_ || _2558_;
  assign _2625_ = _2624_ || _2559_;
  assign _2626_ = _2625_ || _2560_;
  assign _2627_ = _2626_ || _2561_;
  assign _2628_ = _2627_ || _2562_;
  assign _2629_ = _2628_ || _2563_;
  assign _2630_ = _2629_ || _2564_;
  assign _2631_ = _2630_ || _2565_;
  assign _2632_ = _2631_ || _2566_;
  assign _2633_ = _2632_ || _2567_;
  assign _2634_ = _2633_ || _2568_;
  assign _2635_ = _2634_ || _2569_;
  assign _2636_ = _2635_ || _2570_;
  assign _2637_ = _2636_ || _2571_;
  assign _2638_ = _2637_ || _2572_;
  assign _2639_ = _2638_ || _2573_;
  assign _2640_ = _2639_ || _2574_;
  assign _2641_ = _2640_ || _2575_;
  assign _2642_ = _2641_ || _2576_;
  assign _2643_ = _2642_ || _2577_;
  assign _2644_ = _2643_ || _2541_;
  assign _2645_ = _2644_ || _2542_;
  assign _2646_ = _2645_ || _2543_;
  assign _2647_ = _2646_ || _2544_;
  assign _2648_ = _2647_ || _2545_;
  assign _2649_ = _2648_ || _2578_;
  assign _2650_ = _2649_ || _2579_;
  assign _2651_ = _2650_ || _2580_;
  assign _2652_ = _2651_ || _2581_;
  assign _2653_ = _2652_ || _2582_;
  assign \u_frontend.u_decode.u_dec1.rd_valid_o = _2653_ || _2583_;
  assign _2654_ = _2558_ || _2550_;
  assign _2655_ = _2654_ || _2552_;
  assign _2656_ = _2655_ || _2553_;
  assign _2657_ = _2656_ || _2557_;
  assign _2658_ = _2657_ || _2554_;
  assign _2659_ = _2658_ || _2551_;
  assign _2660_ = _2659_ || _2555_;
  assign _2661_ = _2660_ || _2556_;
  assign _2662_ = _2661_ || _2548_;
  assign _2663_ = _2662_ || _2549_;
  assign _2664_ = _2663_ || _2559_;
  assign _2665_ = _2664_ || _2560_;
  assign _2666_ = _2665_ || _2562_;
  assign _2667_ = _2666_ || _2563_;
  assign _2668_ = _2667_ || _2564_;
  assign _2669_ = _2668_ || _2567_;
  assign _2670_ = _2669_ || _2568_;
  assign _2671_ = _2670_ || _2561_;
  assign _2672_ = _2671_ || _2565_;
  assign \u_frontend.u_decode.u_dec1.exec_o = _2672_ || _2566_;
  assign _2673_ = _2569_ || _2570_;
  assign _2674_ = _2673_ || _2571_;
  assign _2675_ = _2674_ || _2572_;
  assign _2676_ = _2675_ || _2573_;
  assign _2677_ = _2676_ || _2574_;
  assign _2678_ = _2677_ || _2584_;
  assign _2679_ = _2678_ || _2585_;
  assign \u_frontend.u_decode.u_dec1.lsu_o = _2679_ || _2586_;
  assign _2680_ = _2613_ || _2587_;
  assign _2681_ = _2680_ || _2588_;
  assign _2682_ = _2681_ || _2589_;
  assign _2683_ = _2682_ || _2590_;
  assign _2684_ = _2683_ || _2591_;
  assign \u_frontend.u_decode.u_dec1.branch_o = _2684_ || _2592_;
  assign _2685_ = _2575_ || _2576_;
  assign _2686_ = _2685_ || _2577_;
  assign _2687_ = _2686_ || _2541_;
  assign _2688_ = _2542_ || _2543_;
  assign _2689_ = _2688_ || _2544_;
  assign _2690_ = _2689_ || _2545_;
  assign _2691_ = _2593_ || _2594_;
  assign _2692_ = _2691_ || _2595_;
  assign _2693_ = _2692_ || _2578_;
  assign _2694_ = _2693_ || _2579_;
  assign _2695_ = _2694_ || _2580_;
  assign _2696_ = _2695_ || _2581_;
  assign _2697_ = _2696_ || _2582_;
  assign _2698_ = _2697_ || _2583_;
  assign _2699_ = _2698_ || _2596_;
  assign _2700_ = _2699_ || _2597_;
  assign _2701_ = _2700_ || _2598_;
  assign _2702_ = _2701_ || _2599_;
  assign _2703_ = _2702_ || \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_frontend.u_decode.u_dec1.csr_o = _2703_ || \u_frontend.u_decode.u_dec1.fetch_fault_i ;
  assign _2704_ = \u_frontend.u_decode.u_dec1.exec_o || _2547_;
  assign _2705_ = _2704_ || _2546_;
  assign _2706_ = _2705_ || _2587_;
  assign _2707_ = _2706_ || _2588_;
  assign _2708_ = _2707_ || _2589_;
  assign _2709_ = _2708_ || _2590_;
  assign _2710_ = _2709_ || _2591_;
  assign _2711_ = _2710_ || _2592_;
  assign _2712_ = _2711_ || _2569_;
  assign _2713_ = _2712_ || _2570_;
  assign _2714_ = _2713_ || _2571_;
  assign _2715_ = _2714_ || _2572_;
  assign _2716_ = _2715_ || _2573_;
  assign _2717_ = _2716_ || _2574_;
  assign _2718_ = _2717_ || _2584_;
  assign _2719_ = _2718_ || _2585_;
  assign _2720_ = _2719_ || _2586_;
  assign _2721_ = _2720_ || _2593_;
  assign _2722_ = _2721_ || _2594_;
  assign _2723_ = _2722_ || _2595_;
  assign _2724_ = _2723_ || _2578_;
  assign _2725_ = _2724_ || _2579_;
  assign _2726_ = _2725_ || _2580_;
  assign _2727_ = _2726_ || _2581_;
  assign _2728_ = _2727_ || _2582_;
  assign _2729_ = _2728_ || _2583_;
  assign _2730_ = _2729_ || _2596_;
  assign _2731_ = _2730_ || _2597_;
  assign _2732_ = _2731_ || _2598_;
  assign _2733_ = _2732_ || _2599_;
  assign _2734_ = _2733_ || _2605_;
  assign _2735_ = _2734_ || _2606_;
  assign _2736_ = _2735_ || _2607_;
  assign _2737_ = ~ _2612_;
  assign _2748_ = \u_frontend.u_decode.u_fifo.wr_ptr_q + 1'h1;
  assign _2749_[0] = \u_frontend.u_decode.u_fifo.rd_ptr_q + 1'h1;
  assign _2750_[1:0] = \u_frontend.u_decode.u_fifo.count_q + 1'h1;
  assign \u_frontend.u_decode.u_fifo.push_w = \u_frontend.u_decode.u_fifo.push_i & \u_frontend.u_decode.u_fifo.accept_o ;
  assign \u_frontend.u_decode.u_fifo.pop1_w = \u_frontend.u_decode.u_fifo.pop0_i & \u_frontend.u_decode.u_dec0.valid_i ;
  assign \u_frontend.u_decode.u_fifo.pop2_w = \u_frontend.u_decode.u_fifo.pop1_i & \u_frontend.u_decode.u_dec1.valid_i ;
  assign _2751_ = \u_frontend.u_decode.u_fifo.push_w & _2762_;
  assign _2752_ = _2763_ & \u_frontend.u_decode.u_fifo.pop_complete_w ;
  assign \u_frontend.u_decode.u_dec0.valid_i = _2759_ & _2757_;
  assign \u_frontend.u_decode.u_dec1.valid_i = _2759_ & _2758_;
  assign _2753_ = \u_frontend.u_decode.u_fifo.pop1_w && _2760_;
  assign _2754_ = \u_frontend.u_decode.u_fifo.pop2_w && _2761_;
  assign _2755_ = \u_frontend.u_decode.u_fifo.pop1_w && \u_frontend.u_decode.u_fifo.pop2_w ;
  assign _2756_ = _2753_ || _2754_;
  assign \u_frontend.u_decode.u_fifo.pop_complete_w = _2756_ || _2755_;
  assign _2759_ = | \u_frontend.u_decode.u_fifo.count_q ;
  assign \u_frontend.u_decode.u_fifo.accept_o = \u_frontend.u_decode.u_fifo.count_q != 2'h2;
  assign _2760_ = ~ \u_frontend.u_decode.u_dec1.valid_i ;
  assign _2761_ = ~ \u_frontend.u_decode.u_dec0.valid_i ;
  assign _2743_ = ~ \u_frontend.u_decode.u_fifo.pred_in_i [0];
  assign _2762_ = ~ \u_frontend.u_decode.u_fifo.pop_complete_w ;
  assign _2763_ = ~ \u_frontend.u_decode.u_fifo.push_w ;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.rd_ptr_q <= _2746_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.wr_ptr_q <= _2747_;
  always @(posedge clk_i)
      \u_frontend.u_decode.u_fifo.count_q <= _2745_;
  assign _2739_[1] = rst_i ? 1'h1 : 1'h0;
  assign _2764_[1] = \u_frontend.u_decode.u_fifo.flush_i ? 1'h1 : 1'h0;
  assign _2740_[1] = rst_i ? 1'h0 : _2764_[1];
  assign _2765_[63] = \u_frontend.u_decode.u_fifo.push_w ? 1'h1 : 1'h0;
  assign _2766_[63] = \u_frontend.u_decode.u_fifo.flush_i ? 1'h0 : _2765_[63];
  assign _2741_[1] = rst_i ? 1'h0 : _2766_[63];
  assign _2767_ = \u_frontend.u_decode.u_fifo.pop1_w ? 1'h1 : 1'h0;
  assign _2768_ = \u_frontend.u_decode.u_fifo.flush_i ? 1'h0 : _2767_;
  assign _2742_ = rst_i ? 1'h0 : _2768_;
  assign _2769_ = \u_frontend.u_decode.u_fifo.pop2_w ? 1'h1 : 1'h0;
  assign _2770_ = \u_frontend.u_decode.u_fifo.flush_i ? 1'h0 : _2769_;
  assign _2744_ = rst_i ? 1'h0 : _2770_;
  assign _2771_ = _2752_ ? _2778_[1:0] : \u_frontend.u_decode.u_fifo.count_q ;
  assign _2772_ = _2751_ ? _2750_[1:0] : _2771_;
  assign _2773_ = \u_frontend.u_decode.u_fifo.flush_i ? 2'h0 : _2772_;
  assign _2745_ = rst_i ? 2'h0 : _2773_;
  assign _2774_ = \u_frontend.u_decode.u_fifo.push_w ? _2748_ : \u_frontend.u_decode.u_fifo.wr_ptr_q ;
  assign _2775_ = \u_frontend.u_decode.u_fifo.flush_i ? 1'h0 : _2774_;
  assign _2747_ = rst_i ? 1'h0 : _2775_;
  assign _2776_ = \u_frontend.u_decode.u_fifo.pop_complete_w ? _2749_[0] : \u_frontend.u_decode.u_fifo.rd_ptr_q ;
  assign _2777_ = \u_frontend.u_decode.u_fifo.flush_i ? 1'h0 : _2776_;
  assign _2746_ = rst_i ? 1'h0 : _2777_;
  assign _2778_[1:0] = \u_frontend.u_decode.u_fifo.count_q - 1'h1;
  assign _2789_ = \u_frontend.u_fetch.branch_q & _2799_;
  assign _2790_ = \u_frontend.u_fetch.branch_w & _2810_;
  assign _2791_ = \u_frontend.u_fetch.active_q & \u_frontend.u_decode.u_fifo.accept_o ;
  assign \u_frontend.u_fetch.icache_rd_o = _2791_ & _2801_;
  assign \u_frontend.u_decode.u_fifo.push_i = _2808_ & _2804_;
  assign _2792_ = \u_frontend.u_decode.u_fifo.flush_i && _2806_;
  assign _2793_ = $signed(32'h00000000) && \u_frontend.u_fetch.branch_w ;
  assign _2794_ = _2793_ && \u_frontend.u_fetch.pc_accept_o ;
  assign _2795_ = \u_frontend.u_fetch.icache_rd_o && mem_i_accept_i;
  assign _2797_ = _2796_ && \u_frontend.u_fetch.branch_w ;
  assign \u_frontend.u_fetch.icache_busy_w = \u_frontend.u_fetch.icache_fetch_q && _2802_;
  assign _2798_ = \u_frontend.u_decode.u_fifo.push_i && _2803_;
  assign _2799_ = ! \u_frontend.u_decode.u_fifo.flush_i ;
  assign _2800_ = ! \u_frontend.u_fetch.active_q ;
  assign _2801_ = ! \u_frontend.u_fetch.icache_busy_w ;
  assign _2802_ = ! mem_i_valid_i;
  assign _2803_ = ! \u_frontend.u_decode.u_fifo.accept_o ;
  assign _2804_ = ! \u_frontend.u_fetch.branch_w ;
  assign _2805_ = ! mem_i_accept_i;
  assign \u_frontend.u_fetch.branch_w = \u_frontend.u_fetch.branch_q || \u_frontend.u_decode.u_fifo.flush_i ;
  assign _2806_ = \u_frontend.u_fetch.icache_busy_w || _2800_;
  assign _2807_ = \u_frontend.u_fetch.stall_w || _2800_;
  assign _2796_ = _2807_ || \u_frontend.u_fetch.stall_q ;
  assign _2808_ = mem_i_valid_i || \u_frontend.u_fetch.skid_valid_q ;
  assign _2809_ = _2803_ || \u_frontend.u_fetch.icache_busy_w ;
  assign \u_frontend.u_fetch.stall_w = _2809_ || _2805_;
  assign \u_frontend.u_fetch.pc_accept_o = ~ \u_frontend.u_fetch.stall_w ;
  assign _2810_ = ~ \u_frontend.u_fetch.stall_q ;
  assign \u_frontend.u_fetch.icache_flush_o = \u_csr.ifence_q | \u_frontend.u_fetch.icache_invalidate_q ;
  always @(posedge clk_i)
      \u_frontend.u_fetch.branch_q <= _2781_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.branch_pc_q <= _2780_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.skid_buffer_q <= _2786_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.skid_valid_q <= _2787_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.pred_d_q <= _2785_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.pc_d_q <= _2783_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.pc_f_q <= _2784_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.icache_invalidate_q <= 1'h0;
  always @(posedge clk_i)
      \u_frontend.u_fetch.icache_fetch_q <= _2782_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.stall_q <= _2788_;
  always @(posedge clk_i)
      \u_frontend.u_fetch.active_q <= _2779_;
  assign _2811_ = \u_frontend.u_fetch.icache_busy_w ? \u_frontend.u_fetch.branch_pc_q : 32'h00000000;
  assign _2812_ = _2792_ ? \u_frontend.u_fetch.branch_pc_w : _2811_;
  assign _2780_ = rst_i ? 32'h00000000 : _2812_;
  assign _2813_ = \u_frontend.u_fetch.icache_busy_w ? \u_frontend.u_fetch.branch_q : 1'h0;
  assign _2814_ = _2792_ ? \u_frontend.u_fetch.branch_w : _2813_;
  assign _2781_ = rst_i ? 1'h0 : _2814_;
  assign _2815_ = _2798_ ? 1'h1 : 1'h0;
  assign _2787_ = rst_i ? 1'h0 : _2815_;
  logic [99:0] fangyuan92;
  assign fangyuan92 = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i , \u_frontend.u_fetch.fetch_pred_branch_o [1], \u_frontend.u_decode.u_fifo.pred_in_i [0], \u_frontend.u_decode.u_fifo.pc_in_i , \u_frontend.u_decode.fetch_in_instr_i };
  assign _2816_ = _2798_ ? fangyuan92 : 100'h0000000000000000000000000;
  assign _2786_ = rst_i ? 100'h0000000000000000000000000 : _2816_;
  assign _2817_ = mem_i_valid_i ? 2'h0 : \u_frontend.u_fetch.pred_d_q ;
  assign _2818_ = _2795_ ? \u_frontend.u_fetch.next_taken_f_i : _2817_;
  assign _2785_ = rst_i ? 2'h0 : _2818_;
  assign _2819_ = _2795_ ? \u_frontend.u_fetch.icache_pc_w : \u_frontend.u_fetch.pc_d_q ;
  assign _2783_ = rst_i ? 32'h00000000 : _2819_;
  assign _2820_ = \u_frontend.u_fetch.stall_w ? \u_frontend.u_fetch.pc_f_q : \u_frontend.u_fetch.next_pc_f_i ;
  assign _2821_ = _2797_ ? \u_frontend.u_fetch.branch_pc_w : _2820_;
  assign _2822_ = _2794_ ? \u_frontend.u_fetch.branch_pc_w : _2821_;
  assign _2784_ = rst_i ? 32'h00000000 : _2822_;
  assign _2823_ = mem_i_valid_i ? 1'h0 : \u_frontend.u_fetch.icache_fetch_q ;
  assign _2824_ = _2795_ ? 1'h1 : _2823_;
  assign _2782_ = rst_i ? 1'h0 : _2824_;
  assign _2788_ = rst_i ? 1'h0 : \u_frontend.u_fetch.stall_w ;
  assign _2825_ = \u_frontend.u_fetch.branch_w ? 1'h1 : \u_frontend.u_fetch.active_q ;
  assign _2826_ = _2794_ ? 1'h1 : _2825_;
  assign _2779_ = rst_i ? 1'h0 : _2826_;
  assign \u_frontend.u_fetch.branch_pc_w = _2789_ ? \u_frontend.u_fetch.branch_pc_q : \u_frontend.u_fetch.branch_pc_i ;
  assign \u_frontend.u_fetch.icache_pc_w = _2790_ ? \u_frontend.u_fetch.branch_pc_w : \u_frontend.u_fetch.pc_f_q ;
  logic [31:0] fangyuan93;
  assign fangyuan93 = { \u_frontend.u_fetch.pc_d_q [31:3], 3'h0 };
  assign \u_frontend.u_decode.u_fifo.pc_in_i = \u_frontend.u_fetch.skid_valid_q ? \u_frontend.u_fetch.skid_buffer_q [95:64] : fangyuan93;
  assign \u_frontend.u_decode.fetch_in_instr_i = \u_frontend.u_fetch.skid_valid_q ? \u_frontend.u_fetch.skid_buffer_q [63:0] : mem_i_inst_i;
  logic [1:0] fangyuan94;
  assign { \u_frontend.u_fetch.fetch_pred_branch_o [1], \u_frontend.u_decode.u_fifo.pred_in_i [0] } = fangyuan94;
  assign fangyuan94 = \u_frontend.u_fetch.skid_valid_q ? \u_frontend.u_fetch.skid_buffer_q [97:96] : \u_frontend.u_fetch.pred_d_q ;
  assign \u_frontend.u_decode.fetch_in_fault_fetch_i = \u_frontend.u_fetch.skid_valid_q ? \u_frontend.u_fetch.skid_buffer_q [98] : mem_i_error_i;
  assign \u_frontend.u_decode.fetch_in_fault_page_i = \u_frontend.u_fetch.skid_valid_q ? \u_frontend.u_fetch.skid_buffer_q [99] : 1'h0;
  assign _2956_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_q + 1'h1;
  assign _2957_[2:0] = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q + 1'h1;
  assign _2835_ = \u_frontend.u_npc.branch_source_i + 3'h4;
  assign _2837_ = _3064_ + 3'h4;
  assign _2828_ = _2999_ + 1'h1;
  logic [31:0] fangyuan95;
  assign fangyuan95 = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign _2958_ = fangyuan95 + 4'h8;
  assign _2959_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r & \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_w ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.ras_call_pred_w = _2959_ & _2966_[0];
  assign _2960_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r & \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_w ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.ras_ret_pred_w = _2960_ & _2966_[0];
  assign _2961_ = \u_frontend.u_npc.branch_request_i & \u_frontend.u_npc.branch_is_call_i ;
  assign _2962_ = \u_frontend.u_npc.branch_request_i & \u_frontend.u_npc.branch_is_ret_i ;
  assign _2963_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_call_pred_w & \u_frontend.u_fetch.pc_accept_o ;
  assign _2964_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_ret_pred_w & \u_frontend.u_fetch.pc_accept_o ;
  assign _2965_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r & _3048_;
  assign _2968_ = _3025_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2969_ = _3026_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2970_ = _3027_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2971_ = _3028_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2972_ = _3029_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2973_ = _3030_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2974_ = _3031_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2975_ = _3032_ == \u_frontend.u_fetch.icache_pc_w ;
  assign _2976_ = _3025_ == _3045_;
  assign _2977_ = _3026_ == _3045_;
  assign _2978_ = _3027_ == _3045_;
  assign _2979_ = _3028_ == _3045_;
  assign _2980_ = _3029_ == _3045_;
  assign _2981_ = _3030_ == _3045_;
  assign _2982_ = _3031_ == _3045_;
  assign _2983_ = _3032_ == _3045_;
  assign _2984_ = _3025_ == \u_frontend.u_npc.branch_source_i ;
  assign _2985_ = _3026_ == \u_frontend.u_npc.branch_source_i ;
  assign _2986_ = _3027_ == \u_frontend.u_npc.branch_source_i ;
  assign _2987_ = _3028_ == \u_frontend.u_npc.branch_source_i ;
  assign _2988_ = _3029_ == \u_frontend.u_npc.branch_source_i ;
  assign _2989_ = _3030_ == \u_frontend.u_npc.branch_source_i ;
  assign _2990_ = _3031_ == \u_frontend.u_npc.branch_source_i ;
  assign _2991_ = _3032_ == \u_frontend.u_npc.branch_source_i ;
  assign _2992_ = _3000_ >= 2'h2;
  assign _2993_ = _2999_ > 1'h0;
  assign _2994_ = \u_frontend.u_npc.branch_is_taken_i && _2998_;
  assign _2995_ = \u_frontend.u_npc.branch_is_not_taken_i && _2993_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.bht_predict_taken_w = $signed(32'h00000001) && _2992_;
  assign _2996_ = _3041_ && _3042_;
  assign _2997_ = _2964_ || _2962_;
  assign _2998_ = _2999_ < 2'h3;
  assign _2966_[0] = ~ \u_frontend.u_npc.BRANCH_PREDICTION.ras_pc_pred_w [0];
  assign _3041_ = ~ _2952_;
  assign _3042_ = ~ \u_frontend.u_fetch.icache_pc_w [2];
  assign _3043_ = ~ _2954_;
  assign _3044_ = ~ \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ;
  assign _3045_ = \u_frontend.u_fetch.icache_pc_w | 3'h4;
  assign _3046_ = \u_frontend.u_npc.BRANCH_PREDICTION.bht_predict_taken_w | \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_r ;
  assign _3047_ = \u_frontend.u_npc.BRANCH_PREDICTION.ras_ret_pred_w | \u_frontend.u_npc.BRANCH_PREDICTION.bht_predict_taken_w ;
  assign _3048_ = _3047_ | \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_r ;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q <= _2839_;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_q <= _2840_;
  assign _2827_[1] = rst_i ? 1'h1 : 1'h0;
  assign _3049_[31] = \u_frontend.u_npc.BRANCH_PREDICTION.btb_hit_r ? 1'h1 : 1'h0;
  assign _2832_ = rst_i ? 1'h0 : _3049_[31];
  assign _3050_[31] = \u_frontend.u_npc.branch_is_taken_i ? 1'h1 : 1'h0;
  assign _3051_[31] = \u_frontend.u_npc.BRANCH_PREDICTION.btb_hit_r ? _3050_[31] : 1'h0;
  assign _2834_[31] = rst_i ? 1'h0 : _3051_[31];
  assign _3052_[31] = \u_frontend.u_npc.BRANCH_PREDICTION.btb_miss_r ? 1'h1 : 1'h0;
  assign _3053_[31] = \u_frontend.u_npc.BRANCH_PREDICTION.btb_hit_r ? 1'h0 : _3052_[31];
  assign _2833_ = rst_i ? 1'h0 : _3053_[31];
  assign _2955_ = _2991_ ? 3'h7 : _2953_;
  assign _2954_ = _2991_ ? 1'h1 : _2946_;
  assign _2953_ = _2990_ ? 3'h6 : _2945_;
  assign _2946_ = _2990_ ? 1'h1 : _2938_;
  assign _2945_ = _2989_ ? 3'h5 : _2937_;
  assign _2938_ = _2989_ ? 1'h1 : _2930_;
  logic [2:0] fangyuan96;
  assign fangyuan96 = { 1'h0, _2929_ };
  assign _2937_ = _2988_ ? 3'h4 : fangyuan96;
  assign _2930_ = _2988_ ? 1'h1 : _2922_;
  assign _2929_ = _2987_ ? 2'h3 : _2920_;
  assign _2922_ = _2987_ ? 1'h1 : _2913_;
  logic [1:0] fangyuan97;
  assign fangyuan97 = { 1'h0, _2911_ };
  assign _2920_ = _2986_ ? 2'h2 : fangyuan97;
  assign _2913_ = _2986_ ? 1'h1 : _2904_;
  assign _2911_ = _2985_ ? 1'h1 : 1'h0;
  assign _2904_ = _2985_ ? 1'h1 : _2895_;
  assign _2895_ = _2984_ ? 1'h1 : 1'h0;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_miss_r = \u_frontend.u_npc.branch_request_i ? _3043_ : 1'h0;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_hit_r = \u_frontend.u_npc.branch_request_i ? _2954_ : 1'h0;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_entry_r = \u_frontend.u_npc.branch_request_i ? _2955_ : 3'h0;
  assign _2886_ = _2983_ ? _3040_ : _2880_;
  assign _2884_ = _2983_ ? _3016_ : _2878_;
  assign _2885_ = _2983_ ? _3024_ : _2879_;
  assign _2883_ = _2983_ ? _3008_ : _2877_;
  assign _2887_ = _2983_ ? 1'h1 : _2881_;
  assign _2888_ = _2983_ ? 1'h1 : _2882_;
  assign _2880_ = _2982_ ? _3039_ : _2874_;
  assign _2878_ = _2982_ ? _3015_ : _2872_;
  assign _2879_ = _2982_ ? _3023_ : _2873_;
  assign _2877_ = _2982_ ? _3007_ : _2871_;
  assign _2881_ = _2982_ ? 1'h1 : _2875_;
  assign _2882_ = _2982_ ? 1'h1 : _2876_;
  assign _2874_ = _2981_ ? _3038_ : _2868_;
  assign _2872_ = _2981_ ? _3014_ : _2866_;
  assign _2873_ = _2981_ ? _3022_ : _2867_;
  assign _2871_ = _2981_ ? _3006_ : _2865_;
  assign _2875_ = _2981_ ? 1'h1 : _2869_;
  assign _2876_ = _2981_ ? 1'h1 : _2870_;
  assign _2868_ = _2980_ ? _3037_ : _2862_;
  assign _2866_ = _2980_ ? _3013_ : _2860_;
  assign _2867_ = _2980_ ? _3021_ : _2861_;
  assign _2865_ = _2980_ ? _3005_ : _2859_;
  assign _2869_ = _2980_ ? 1'h1 : _2863_;
  assign _2870_ = _2980_ ? 1'h1 : _2864_;
  assign _2862_ = _2979_ ? _3036_ : _2856_;
  assign _2860_ = _2979_ ? _3012_ : _2854_;
  assign _2861_ = _2979_ ? _3020_ : _2855_;
  assign _2859_ = _2979_ ? _3004_ : _2853_;
  assign _2863_ = _2979_ ? 1'h1 : _2857_;
  assign _2864_ = _2979_ ? 1'h1 : _2858_;
  assign _2856_ = _2978_ ? _3035_ : _2850_;
  assign _2854_ = _2978_ ? _3011_ : _2848_;
  assign _2855_ = _2978_ ? _3019_ : _2849_;
  assign _2853_ = _2978_ ? _3003_ : _2847_;
  assign _2857_ = _2978_ ? 1'h1 : _2851_;
  assign _2858_ = _2978_ ? 1'h1 : _2852_;
  assign _2850_ = _2977_ ? _3034_ : _2844_;
  assign _2848_ = _2977_ ? _3010_ : _2842_;
  assign _2849_ = _2977_ ? _3018_ : _2843_;
  assign _2847_ = _2977_ ? _3002_ : _2841_;
  assign _2851_ = _2977_ ? 1'h1 : _2845_;
  assign _2852_ = _2977_ ? 1'h1 : _2846_;
  assign _2844_ = _2976_ ? _3033_ : _2950_;
  assign _2842_ = _2976_ ? _3009_ : _2948_;
  assign _2843_ = _2976_ ? _3017_ : _2949_;
  assign _2841_ = _2976_ ? _3001_ : _2947_;
  assign _2845_ = _2976_ ? 1'h1 : _2951_;
  assign _2846_ = _2976_ ? 1'h1 : _2952_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_jmp_r = _2996_ ? _2884_ : _2948_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_next_pc_r = _2996_ ? _2886_ : _2950_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_w = _2996_ ? _2885_ : _2949_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_w = _2996_ ? _2883_ : _2947_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r = _2996_ ? _2887_ : _2951_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r = _2996_ ? _2888_ : _2952_;
  assign _2950_ = _2975_ ? _3040_ : _2942_;
  assign _2948_ = _2975_ ? _3016_ : _2940_;
  assign _2949_ = _2975_ ? _3024_ : _2941_;
  assign _2947_ = _2975_ ? _3008_ : _2939_;
  assign _2951_ = _2975_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2943_;
  assign _2952_ = _2975_ ? 1'h1 : _2944_;
  assign _2942_ = _2974_ ? _3039_ : _2934_;
  assign _2940_ = _2974_ ? _3015_ : _2932_;
  assign _2941_ = _2974_ ? _3023_ : _2933_;
  assign _2939_ = _2974_ ? _3007_ : _2931_;
  assign _2943_ = _2974_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2935_;
  assign _2944_ = _2974_ ? 1'h1 : _2936_;
  assign _2934_ = _2973_ ? _3038_ : _2926_;
  assign _2932_ = _2973_ ? _3014_ : _2924_;
  assign _2933_ = _2973_ ? _3022_ : _2925_;
  assign _2931_ = _2973_ ? _3006_ : _2923_;
  assign _2935_ = _2973_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2927_;
  assign _2936_ = _2973_ ? 1'h1 : _2928_;
  assign _2926_ = _2972_ ? _3037_ : _2917_;
  assign _2924_ = _2972_ ? _3013_ : _2915_;
  assign _2925_ = _2972_ ? _3021_ : _2916_;
  assign _2923_ = _2972_ ? _3005_ : _2914_;
  assign _2927_ = _2972_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2918_;
  assign _2928_ = _2972_ ? 1'h1 : _2919_;
  assign _2917_ = _2971_ ? _3036_ : _2908_;
  assign _2915_ = _2971_ ? _3012_ : _2906_;
  assign _2916_ = _2971_ ? _3020_ : _2907_;
  assign _2914_ = _2971_ ? _3004_ : _2905_;
  assign _2918_ = _2971_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2909_;
  assign _2919_ = _2971_ ? 1'h1 : _2910_;
  assign _2908_ = _2970_ ? _3035_ : _2899_;
  assign _2906_ = _2970_ ? _3011_ : _2897_;
  assign _2907_ = _2970_ ? _3019_ : _2898_;
  assign _2905_ = _2970_ ? _3003_ : _2896_;
  assign _2909_ = _2970_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2900_;
  assign _2910_ = _2970_ ? 1'h1 : _2901_;
  assign _2899_ = _2969_ ? _3034_ : _2892_;
  assign _2897_ = _2969_ ? _3010_ : _2890_;
  assign _2898_ = _2969_ ? _3018_ : _2891_;
  assign _2896_ = _2969_ ? _3002_ : _2889_;
  assign _2900_ = _2969_ ? \u_frontend.u_fetch.icache_pc_w [2] : _2893_;
  assign _2901_ = _2969_ ? 1'h1 : _2894_;
  assign _2892_ = _2968_ ? _3033_ : _2958_;
  assign _2890_ = _2968_ ? _3009_ : 1'h0;
  assign _2891_ = _2968_ ? _3017_ : 1'h0;
  assign _2889_ = _2968_ ? _3001_ : 1'h0;
  assign _2893_ = _2968_ ? \u_frontend.u_fetch.icache_pc_w [2] : 1'h0;
  assign _2894_ = _2968_ ? 1'h1 : 1'h0;
  assign _3054_[1] = _2994_ ? 1'h1 : 1'h0;
  assign _2829_[1] = rst_i ? 1'h0 : _3054_[1];
  assign _3055_[1] = _2995_ ? 1'h1 : 1'h0;
  assign _3056_[1] = _2994_ ? 1'h0 : _3055_[1];
  assign _2831_[1] = rst_i ? 1'h0 : _3056_[1];
  assign _3057_[31] = _2961_ ? 1'h1 : 1'h0;
  assign _2836_[31] = rst_i ? 1'h0 : _3057_[31];
  assign _3058_[31] = _2963_ ? 1'h1 : 1'h0;
  assign _3059_[31] = _2961_ ? 1'h0 : _3058_[31];
  assign _2838_[31] = rst_i ? 1'h0 : _3059_[31];
  assign _3060_ = _2997_ ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r : \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q ;
  assign _3061_ = _2963_ ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r : _3060_;
  assign _3062_ = _2961_ ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r : _3061_;
  assign _2839_ = rst_i ? 3'h0 : _3062_;
  assign _2921_ = _2964_ ? _3063_[2:0] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q ;
  assign _2912_ = _2963_ ? _2957_[2:0] : _2921_;
  assign _2902_ = _2962_ ? _2967_[2:0] : _2912_;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_r = _2961_ ? _2956_ : _2902_;
  assign _2840_ = rst_i ? 3'h0 : \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_r ;
  assign _2903_ = _2962_ ? _2967_[2:0] : \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_q ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_r = _2961_ ? _2956_ : _2903_;
  assign _2967_[2:0] = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_real_q - 1'h1;
  assign _3063_[2:0] = \u_frontend.u_npc.BRANCH_PREDICTION.ras_index_q - 1'h1;
  assign _2830_ = _2999_ - 1'h1;
  assign _3064_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ? _3045_ : \u_frontend.u_fetch.icache_pc_w ;
  assign _3065_ = _3046_ ? \u_frontend.u_npc.BRANCH_PREDICTION.btb_next_pc_r : _2958_;
  assign \u_frontend.u_fetch.next_pc_f_i = \u_frontend.u_npc.BRANCH_PREDICTION.ras_ret_pred_w ? \u_frontend.u_npc.BRANCH_PREDICTION.ras_pc_pred_w : _3065_;
  assign _3066_[0] = \u_frontend.u_fetch.icache_pc_w [2] ? 1'h0 : _3044_;
  logic [1:0] fangyuan98;
  assign fangyuan98 = { \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r , _3066_[0] };
  assign \u_frontend.u_fetch.next_taken_f_i = _2965_ ? fangyuan98 : 2'h0;
  always @(posedge clk_i)
      \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q <= _3067_;
  logic [15:0] fangyuan99;
  assign fangyuan99 = { 1'h0, \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [15:1] };
  assign _3068_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [0] ? _3070_ : fangyuan99;
  assign _3069_ = \u_frontend.u_npc.BRANCH_PREDICTION.btb_miss_r ? _3068_ : \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q ;
  assign _3067_ = rst_i ? 16'h0001 : _3069_;
  assign _3070_ = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [15:1] ^ 16'hb400;
  assign _3121_ = \u_issue.pc_x_q + 4'h8;
  assign _3122_ = \u_issue.pc_x_q + 3'h4;
  assign _3123_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_taken_q ;
  assign _3124_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] & \u_exec0.branch_taken_q ;
  assign _3125_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_ntaken_q ;
  assign _3126_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] & \u_exec0.branch_ntaken_q ;
  assign _3127_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_call_q ;
  assign _3128_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] & \u_exec0.branch_call_q ;
  assign _3129_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_ret_q ;
  assign _3130_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] & \u_exec0.branch_ret_q ;
  assign _3131_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_jmp_q ;
  assign _3132_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] & \u_exec0.branch_jmp_q ;
  assign _3133_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] & \u_exec1.branch_request_o ;
  assign \u_issue.lsu_opcode_valid_o = _3425_ & _3301_;
  assign \u_issue.dual_issue_w = \u_exec1.opcode_valid_i & _3301_;
  assign _3134_ = \u_div.opcode_valid_i & _3302_;
  assign \u_issue.single_issue_w = _3134_ & _3301_;
  assign _3135_ = \u_issue.slot0_valid_r & \u_div.opcode_valid_i ;
  assign \u_frontend.u_decode.u_fifo.pop0_i = _3308_ & _3301_;
  assign _3136_ = \u_issue.slot1_valid_r & \u_div.opcode_valid_i ;
  assign \u_frontend.u_decode.u_fifo.pop1_i = _3309_ & _3301_;
  assign \u_csr.opcode_valid_i = \u_div.opcode_valid_i & _3301_;
  logic [30:0] fangyuan100;
  assign fangyuan100 = { _3341_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3137_ = | fangyuan100;
  logic [30:0] fangyuan101;
  assign fangyuan101 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3345_, _3344_, _3343_, _3342_ };
  assign _3138_ = | fangyuan101;
  logic [30:0] fangyuan102;
  assign fangyuan102 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3313_, _3312_, _3311_, _3310_ };
  assign _3139_ = | fangyuan102;
  logic [30:0] fangyuan103;
  assign fangyuan103 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3140_ = | fangyuan103;
  logic [30:0] fangyuan104;
  assign fangyuan104 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3141_ = | fangyuan104;
  logic [30:0] fangyuan105;
  assign fangyuan105 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3142_ = | fangyuan105;
  logic [30:0] fangyuan106;
  assign fangyuan106 = { _3373_, _3372_, _3371_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3143_ = | fangyuan106;
  logic [30:0] fangyuan107;
  assign fangyuan107 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3144_ = | fangyuan107;
  logic [30:0] fangyuan108;
  assign fangyuan108 = { _3405_, _3404_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3145_ = | fangyuan108;
  logic [30:0] fangyuan109;
  assign fangyuan109 = { _3341_, _3340_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3146_ = | fangyuan109;
  logic [30:0] fangyuan110;
  assign fangyuan110 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3147_ = | fangyuan110;
  logic [30:0] fangyuan111;
  assign fangyuan111 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3148_ = | fangyuan111;
  logic [30:0] fangyuan112;
  assign fangyuan112 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3149_ = | fangyuan112;
  logic [30:0] fangyuan113;
  assign fangyuan113 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3150_ = | fangyuan113;
  logic [30:0] fangyuan114;
  assign fangyuan114 = { _3373_, _3372_, _3371_, _3370_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3151_ = | fangyuan114;
  logic [30:0] fangyuan115;
  assign fangyuan115 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3152_ = | fangyuan115;
  logic [30:0] fangyuan116;
  assign fangyuan116 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3376_, _3375_, _3374_ };
  assign _3153_ = | fangyuan116;
  logic [30:0] fangyuan117;
  assign fangyuan117 = { _3373_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3154_ = | fangyuan117;
  logic [30:0] fangyuan118;
  assign fangyuan118 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3155_ = | fangyuan118;
  logic [30:0] fangyuan119;
  assign fangyuan119 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3156_ = | fangyuan119;
  logic [30:0] fangyuan120;
  assign fangyuan120 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3157_ = | fangyuan120;
  logic [30:0] fangyuan121;
  assign fangyuan121 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3158_ = | fangyuan121;
  logic [30:0] fangyuan122;
  assign fangyuan122 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3159_ = | fangyuan122;
  logic [30:0] fangyuan123;
  assign fangyuan123 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3160_ = | fangyuan123;
  logic [30:0] fangyuan124;
  assign fangyuan124 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3161_ = | fangyuan124;
  logic [30:0] fangyuan125;
  assign fangyuan125 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3162_ = | fangyuan125;
  logic [30:0] fangyuan126;
  assign fangyuan126 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3163_ = | fangyuan126;
  logic [30:0] fangyuan127;
  assign fangyuan127 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3164_ = | fangyuan127;
  logic [30:0] fangyuan128;
  assign fangyuan128 = { _3373_, _3372_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3165_ = | fangyuan128;
  logic [30:0] fangyuan129;
  assign fangyuan129 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3166_ = | fangyuan129;
  logic [30:0] fangyuan130;
  assign fangyuan130 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_ };
  assign _3167_ = | fangyuan130;
  logic [30:0] fangyuan131;
  assign fangyuan131 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3168_ = | fangyuan131;
  logic [30:0] fangyuan132;
  assign fangyuan132 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3169_ = | fangyuan132;
  logic [30:0] fangyuan133;
  assign fangyuan133 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3170_ = | fangyuan133;
  logic [30:0] fangyuan134;
  assign fangyuan134 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3171_ = | fangyuan134;
  logic [30:0] fangyuan135;
  assign fangyuan135 = { _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3172_ = | fangyuan135;
  logic [30:0] fangyuan136;
  assign fangyuan136 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3173_ = | fangyuan136;
  logic [30:0] fangyuan137;
  assign fangyuan137 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3174_ = | fangyuan137;
  logic [30:0] fangyuan138;
  assign fangyuan138 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3342_ };
  assign _3175_ = | fangyuan138;
  logic [30:0] fangyuan139;
  assign fangyuan139 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3176_ = | fangyuan139;
  logic [30:0] fangyuan140;
  assign fangyuan140 = { _3341_, _3340_, _3339_, _3338_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3177_ = | fangyuan140;
  logic [30:0] fangyuan141;
  assign fangyuan141 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3178_ = | fangyuan141;
  logic [30:0] fangyuan142;
  assign fangyuan142 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3179_ = | fangyuan142;
  logic [30:0] fangyuan143;
  assign fangyuan143 = { _3405_, _3404_, _3403_, _3402_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3180_ = | fangyuan143;
  logic [30:0] fangyuan144;
  assign fangyuan144 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3181_ = | fangyuan144;
  logic [30:0] fangyuan145;
  assign fangyuan145 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3182_ = | fangyuan145;
  logic [30:0] fangyuan146;
  assign fangyuan146 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3183_ = | fangyuan146;
  logic [30:0] fangyuan147;
  assign fangyuan147 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3184_ = | fangyuan147;
  logic [30:0] fangyuan148;
  assign fangyuan148 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3185_ = | fangyuan148;
  logic [30:0] fangyuan149;
  assign fangyuan149 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3186_ = | fangyuan149;
  logic [30:0] fangyuan150;
  assign fangyuan150 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3187_ = | fangyuan150;
  logic [30:0] fangyuan151;
  assign fangyuan151 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3310_ };
  assign _3188_ = | fangyuan151;
  logic [30:0] fangyuan152;
  assign fangyuan152 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3189_ = | fangyuan152;
  logic [30:0] fangyuan153;
  assign fangyuan153 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3344_, _3343_, _3342_ };
  assign _3190_ = | fangyuan153;
  logic [30:0] fangyuan154;
  assign fangyuan154 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3191_ = | fangyuan154;
  logic [30:0] fangyuan155;
  assign fangyuan155 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3192_ = | fangyuan155;
  logic [30:0] fangyuan156;
  assign fangyuan156 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3193_ = | fangyuan156;
  logic [30:0] fangyuan157;
  assign fangyuan157 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3194_ = | fangyuan157;
  logic [30:0] fangyuan158;
  assign fangyuan158 = { _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3195_ = | fangyuan158;
  logic [30:0] fangyuan159;
  assign fangyuan159 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3196_ = | fangyuan159;
  logic [30:0] fangyuan160;
  assign fangyuan160 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3197_ = | fangyuan160;
  logic [30:0] fangyuan161;
  assign fangyuan161 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3198_ = | fangyuan161;
  logic [30:0] fangyuan162;
  assign fangyuan162 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3199_ = | fangyuan162;
  logic [30:0] fangyuan163;
  assign fangyuan163 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3200_ = | fangyuan163;
  logic [30:0] fangyuan164;
  assign fangyuan164 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3201_ = | fangyuan164;
  logic [30:0] fangyuan165;
  assign fangyuan165 = { _3405_, _3404_, _3403_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3202_ = | fangyuan165;
  logic [30:0] fangyuan166;
  assign fangyuan166 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3203_ = | fangyuan166;
  logic [30:0] fangyuan167;
  assign fangyuan167 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3343_, _3342_ };
  assign _3204_ = | fangyuan167;
  logic [30:0] fangyuan168;
  assign fangyuan168 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3374_ };
  assign _3205_ = | fangyuan168;
  logic [30:0] fangyuan169;
  assign fangyuan169 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3206_ = | fangyuan169;
  logic [30:0] fangyuan170;
  assign fangyuan170 = { _3405_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3207_ = | fangyuan170;
  logic [30:0] fangyuan171;
  assign fangyuan171 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3208_ = | fangyuan171;
  logic [30:0] fangyuan172;
  assign fangyuan172 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3375_, _3374_ };
  assign _3209_ = | fangyuan172;
  logic [30:0] fangyuan173;
  assign fangyuan173 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3210_ = | fangyuan173;
  logic [30:0] fangyuan174;
  assign fangyuan174 = { _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3211_ = | fangyuan174;
  logic [30:0] fangyuan175;
  assign fangyuan175 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3212_ = | fangyuan175;
  logic [30:0] fangyuan176;
  assign fangyuan176 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3213_ = | fangyuan176;
  logic [30:0] fangyuan177;
  assign fangyuan177 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_ };
  assign _3214_ = | fangyuan177;
  logic [30:0] fangyuan178;
  assign fangyuan178 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3215_ = | fangyuan178;
  logic [30:0] fangyuan179;
  assign fangyuan179 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3311_, _3310_ };
  assign _3216_ = | fangyuan179;
  logic [30:0] fangyuan180;
  assign fangyuan180 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3217_ = | fangyuan180;
  logic [30:0] fangyuan181;
  assign fangyuan181 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3218_ = | fangyuan181;
  logic [30:0] fangyuan182;
  assign fangyuan182 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3377_, _3376_, _3375_, _3374_ };
  assign _3219_ = | fangyuan182;
  logic [30:0] fangyuan183;
  assign fangyuan183 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3220_ = | fangyuan183;
  logic [30:0] fangyuan184;
  assign fangyuan184 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3221_ = | fangyuan184;
  logic [30:0] fangyuan185;
  assign fangyuan185 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3222_ = | fangyuan185;
  logic [30:0] fangyuan186;
  assign fangyuan186 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3223_ = | fangyuan186;
  logic [30:0] fangyuan187;
  assign fangyuan187 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3224_ = | fangyuan187;
  logic [30:0] fangyuan188;
  assign fangyuan188 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3225_ = | fangyuan188;
  logic [30:0] fangyuan189;
  assign fangyuan189 = { _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_, _3354_, _3353_, _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_ };
  assign _3226_ = | fangyuan189;
  logic [30:0] fangyuan190;
  assign fangyuan190 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_ };
  assign _3227_ = | fangyuan190;
  logic [30:0] fangyuan191;
  assign fangyuan191 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3228_ = | fangyuan191;
  logic [30:0] fangyuan192;
  assign fangyuan192 = { _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_ };
  assign _3229_ = | fangyuan192;
  logic [30:0] fangyuan193;
  assign fangyuan193 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3230_ = | fangyuan193;
  logic [30:0] fangyuan194;
  assign fangyuan194 = { _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3312_, _3311_, _3310_ };
  assign _3231_ = | fangyuan194;
  logic [30:0] fangyuan195;
  assign fangyuan195 = { _3341_, _3340_, _3339_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_ };
  assign _3232_ = | fangyuan195;
  logic [29:0] fangyuan196;
  assign fangyuan196 = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 1'h0 };
  assign _3235_ = fangyuan196 == \u_issue.pc_x_q [31:2];
  logic [29:0] fangyuan197;
  assign fangyuan197 = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 1'h1 };
  assign _3236_ = fangyuan197 == \u_issue.pc_x_q [31:2];
  assign _3237_ = \u_issue.pipe0_rd_wb_w == \u_csr.opcode_opcode_i [19:15];
  assign _3238_ = \u_issue.pipe0_rd_wb_w == \u_csr.opcode_opcode_i [24:20];
  assign _3239_ = \u_issue.pipe1_rd_wb_w == \u_csr.opcode_opcode_i [19:15];
  assign _3240_ = \u_issue.pipe1_rd_wb_w == \u_csr.opcode_opcode_i [24:20];
  assign _3241_ = \u_issue.pipe0_rd_e2_w == \u_csr.opcode_opcode_i [19:15];
  assign _3242_ = \u_issue.pipe0_rd_e2_w == \u_csr.opcode_opcode_i [24:20];
  assign _3243_ = \u_issue.pipe1_rd_e2_w == \u_csr.opcode_opcode_i [19:15];
  assign _3244_ = \u_issue.pipe1_rd_e2_w == \u_csr.opcode_opcode_i [24:20];
  assign _3245_ = \u_issue.pipe0_rd_e1_w == \u_csr.opcode_opcode_i [19:15];
  assign _3246_ = \u_issue.pipe0_rd_e1_w == \u_csr.opcode_opcode_i [24:20];
  assign _3247_ = \u_issue.pipe1_rd_e1_w == \u_csr.opcode_opcode_i [19:15];
  assign _3248_ = \u_issue.pipe1_rd_e1_w == \u_csr.opcode_opcode_i [24:20];
  assign _3249_ = ! \u_csr.opcode_opcode_i [19:15];
  assign _3250_ = ! \u_csr.opcode_opcode_i [24:20];
  assign _3251_ = \u_issue.pipe0_rd_wb_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3252_ = \u_issue.pipe0_rd_wb_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3253_ = \u_issue.pipe1_rd_wb_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3254_ = \u_issue.pipe1_rd_wb_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3255_ = \u_issue.pipe0_rd_e2_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3256_ = \u_issue.pipe0_rd_e2_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3257_ = \u_issue.pipe1_rd_e2_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3258_ = \u_issue.pipe1_rd_e2_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3259_ = \u_issue.pipe0_rd_e1_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3260_ = \u_issue.pipe0_rd_e1_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3261_ = \u_issue.pipe1_rd_e1_w == \u_exec1.opcode_opcode_i [19:15];
  assign _3262_ = \u_issue.pipe1_rd_e1_w == \u_exec1.opcode_opcode_i [24:20];
  assign _3263_ = ! \u_exec1.opcode_opcode_i [19:15];
  assign _3264_ = ! \u_exec1.opcode_opcode_i [24:20];
  assign _3265_ = \u_frontend.u_decode.u_dec0.valid_i && _3235_;
  assign _3266_ = \u_frontend.u_decode.u_dec1.valid_i && _3236_;
  assign _3267_ = \u_div.opcode_valid_i && \u_issue.issue_a_div_w ;
  assign _3268_ = \u_csr.opcode_valid_i && \u_issue.issue_a_csr_w ;
  assign _3269_ = _3306_ && \u_frontend.u_decode.u_dec1.exec_o ;
  assign _3270_ = _3306_ && \u_frontend.u_decode.u_dec1.branch_o ;
  assign _3271_ = _3307_ && \u_frontend.u_decode.u_dec1.lsu_o ;
  assign _3272_ = _3305_ && \u_frontend.u_decode.u_dec1.mul_o ;
  assign _3273_ = \u_issue.pipe1_ok_w && _3286_;
  assign \u_issue.dual_issue_ok_w = _3273_ && _3301_;
  assign _3274_ = _3291_ && _3293_;
  assign _3275_ = \u_issue.opcode_a_valid_r && _3280_;
  assign _3276_ = \u_issue.issue_a_sb_alloc_w && _3418_;
  assign _3277_ = \u_issue.dual_issue_ok_w && \u_issue.opcode_b_valid_r ;
  assign _3278_ = _3277_ && \u_div.opcode_valid_i ;
  assign _3279_ = _3278_ && _3281_;
  assign \u_csr.opcode_invalid_i = \u_div.opcode_valid_i && \u_issue.issue_a_invalid_w ;
  assign _3280_ = ! _3298_;
  assign _3281_ = ! _3300_;
  assign _3282_ = \u_csr.branch_q || \u_issue.squash_w ;
  assign _3283_ = \u_frontend.u_decode.u_dec0.valid_i || \u_frontend.u_decode.u_dec1.valid_i ;
  assign \u_issue.squash_w = \u_issue.pipe0_squash_e1_e2_w || \u_issue.pipe1_squash_e1_e2_w ;
  assign _3284_ = _3269_ || _3270_;
  assign _3285_ = _3284_ || _3271_;
  assign _3286_ = _3285_ || _3272_;
  assign _3287_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [1] || \u_issue.u_pipe0_ctrl.ctrl_e1_q [5];
  assign _3288_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [1] || \u_issue.u_pipe1_ctrl.ctrl_e1_q [5];
  assign _3289_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [1] || \u_issue.u_pipe0_ctrl.ctrl_e1_q [2];
  assign _3290_ = _3289_ || \u_issue.u_pipe1_ctrl.ctrl_e1_q [1];
  assign _3291_ = _3290_ || \u_issue.u_pipe1_ctrl.ctrl_e1_q [2];
  assign _3292_ = \u_issue.issue_a_mul_w || \u_issue.issue_a_div_w ;
  assign _3293_ = _3292_ || \u_issue.issue_a_csr_w ;
  assign _3294_ = \u_issue.lsu_stall_i || \u_exec0.hold_i ;
  assign _3295_ = _3294_ || \u_issue.div_pending_q ;
  assign _3296_ = _3295_ || \u_issue.csr_pending_q ;
  assign _3297_ = _3419_ || _3420_;
  assign _3298_ = _3297_ || _3421_;
  assign _3299_ = _3422_ || _3423_;
  assign _3300_ = _3299_ || _3424_;
  assign \u_csr.interrupt_inhibit_i = \u_issue.csr_pending_q || \u_issue.issue_a_csr_w ;
  assign _3301_ = ~ \u_csr.take_interrupt_q ;
  assign _3302_ = ~ \u_issue.dual_issue_w ;
  assign \u_frontend.u_decode.u_fifo.flush_i = \u_csr.branch_q | \u_frontend.u_npc.branch_request_i ;
  assign \u_csr.u_csrfile.exception_i = \u_issue.u_pipe0_ctrl.exception_wb_q | \u_issue.u_pipe1_ctrl.exception_wb_q ;
  assign \u_frontend.u_npc.branch_is_taken_i = _3123_ | _3124_;
  assign \u_frontend.u_npc.branch_is_not_taken_i = _3125_ | _3126_;
  assign \u_frontend.u_npc.branch_is_call_i = _3127_ | _3128_;
  assign \u_frontend.u_npc.branch_is_ret_i = _3129_ | _3130_;
  assign \u_frontend.u_npc.branch_is_jmp_i = _3131_ | _3132_;
  assign _3303_ = \u_frontend.u_decode.u_dec1.exec_o | \u_frontend.u_decode.u_dec1.branch_o ;
  assign _3304_ = _3303_ | \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_issue.pipe1_ok_w = _3304_ | \u_frontend.u_decode.u_dec1.mul_o ;
  assign _3305_ = \u_issue.issue_a_exec_w | \u_issue.issue_a_lsu_w ;
  assign _3306_ = _3305_ | \u_issue.issue_a_mul_w ;
  assign _3307_ = \u_issue.issue_a_exec_w | \u_issue.issue_a_mul_w ;
  assign _3308_ = _3135_ | \u_issue.slot1_valid_r ;
  assign _3309_ = _3136_ | \u_exec1.opcode_valid_i ;
  assign \u_exec0.hold_i = \u_issue.pipe0_stall_raw_w | \u_issue.pipe1_stall_raw_w ;
  always @(posedge clk_i)
      \u_issue.csr_pending_q <= _3071_;
  always @(posedge clk_i)
      \u_issue.div_pending_q <= _3072_;
  always @(posedge clk_i)
      \u_issue.pc_x_q <= _3073_;
  assign \u_exec1.opcode_rb_operand_i = _3264_ ? 32'h00000000 : _3116_;
  assign \u_exec1.opcode_ra_operand_i = _3263_ ? 32'h00000000 : _3115_;
  assign _3116_ = _3262_ ? \u_exec1.result_q : _3111_;
  assign _3115_ = _3261_ ? \u_exec1.result_q : _3110_;
  assign _3111_ = _3260_ ? \u_exec0.result_q : _3105_;
  assign _3110_ = _3259_ ? \u_exec0.result_q : _3104_;
  assign _3105_ = _3258_ ? \u_issue.pipe1_result_e2_w : _3098_;
  assign _3104_ = _3257_ ? \u_issue.pipe1_result_e2_w : _3097_;
  assign _3098_ = _3256_ ? \u_issue.pipe0_result_e2_w : _3082_;
  assign _3097_ = _3255_ ? \u_issue.pipe0_result_e2_w : _3081_;
  assign _3082_ = _3254_ ? \u_issue.u_pipe1_ctrl.result_wb_q : _3077_;
  assign _3081_ = _3253_ ? \u_issue.u_pipe1_ctrl.result_wb_q : _3076_;
  assign _3077_ = _3252_ ? \u_issue.u_pipe0_ctrl.result_wb_q : \u_issue.issue_b_rb_value_w ;
  assign _3076_ = _3251_ ? \u_issue.u_pipe0_ctrl.result_wb_q : \u_issue.issue_b_ra_value_w ;
  assign \u_div.opcode_rb_operand_i = _3250_ ? 32'h00000000 : _3114_;
  assign \u_csr.opcode_ra_operand_i = _3249_ ? 32'h00000000 : _3113_;
  assign _3114_ = _3248_ ? \u_exec1.result_q : _3109_;
  assign _3113_ = _3247_ ? \u_exec1.result_q : _3108_;
  assign _3109_ = _3246_ ? \u_exec0.result_q : _3103_;
  assign _3108_ = _3245_ ? \u_exec0.result_q : _3102_;
  assign _3103_ = _3244_ ? \u_issue.pipe1_result_e2_w : _3096_;
  assign _3102_ = _3243_ ? \u_issue.pipe1_result_e2_w : _3095_;
  assign _3096_ = _3242_ ? \u_issue.pipe0_result_e2_w : _3080_;
  assign _3095_ = _3241_ ? \u_issue.pipe0_result_e2_w : _3079_;
  assign _3080_ = _3240_ ? \u_issue.u_pipe1_ctrl.result_wb_q : _3075_;
  assign _3079_ = _3239_ ? \u_issue.u_pipe1_ctrl.result_wb_q : _3074_;
  assign _3075_ = _3238_ ? \u_issue.u_pipe0_ctrl.result_wb_q : \u_issue.issue_a_rb_value_w ;
  assign _3074_ = _3237_ ? \u_issue.u_pipe0_ctrl.result_wb_q : \u_issue.issue_a_ra_value_w ;
  assign _3091_ = _3279_ ? \u_frontend.u_decode.u_dec1.mul_o : 1'h0;
  assign _3090_ = _3279_ ? \u_frontend.u_decode.u_dec1.lsu_o : 1'h0;
  assign _3089_ = _3279_ ? 1'h1 : 1'h0;
  assign \u_issue.pipe1_mux_mul_r = _3296_ ? 1'h0 : _3091_;
  assign \u_issue.pipe1_mux_lsu_r = _3296_ ? 1'h0 : _3090_;
  assign \u_exec1.opcode_valid_i = _3296_ ? 1'h0 : _3089_;
  logic [1:0] fangyuan198;
  assign fangyuan198 = { 1'h1, _3112_[30] };
  logic [1:0] fangyuan199;
  assign fangyuan199 = { _3311_, _3188_ };
  always @(1'hx or fangyuan198 or fangyuan199) begin
    casez (fangyuan199)
      2'b?1 :
        _3120_[30] = fangyuan198 [0:0] ;
      2'b1? :
        _3120_[30] = fangyuan198 [1:1] ;
      default:
        _3120_[30] = 1'hx ;
    endcase
  end
  assign _3310_ = \u_csr.opcode_opcode_i [11:7] == 5'h1f;
  assign _3311_ = \u_csr.opcode_opcode_i [11:7] == 5'h1e;
  assign _3312_ = \u_csr.opcode_opcode_i [11:7] == 5'h1d;
  assign _3313_ = \u_csr.opcode_opcode_i [11:7] == 5'h1c;
  assign _3314_ = \u_csr.opcode_opcode_i [11:7] == 5'h1b;
  assign _3315_ = \u_csr.opcode_opcode_i [11:7] == 5'h1a;
  assign _3316_ = \u_csr.opcode_opcode_i [11:7] == 5'h19;
  assign _3317_ = \u_csr.opcode_opcode_i [11:7] == 5'h18;
  assign _3318_ = \u_csr.opcode_opcode_i [11:7] == 5'h17;
  assign _3319_ = \u_csr.opcode_opcode_i [11:7] == 5'h16;
  assign _3320_ = \u_csr.opcode_opcode_i [11:7] == 5'h15;
  assign _3321_ = \u_csr.opcode_opcode_i [11:7] == 5'h14;
  assign _3322_ = \u_csr.opcode_opcode_i [11:7] == 5'h13;
  assign _3323_ = \u_csr.opcode_opcode_i [11:7] == 5'h12;
  assign _3324_ = \u_csr.opcode_opcode_i [11:7] == 5'h11;
  assign _3325_ = \u_csr.opcode_opcode_i [11:7] == 5'h10;
  assign _3326_ = \u_csr.opcode_opcode_i [11:7] == 4'hf;
  assign _3327_ = \u_csr.opcode_opcode_i [11:7] == 4'he;
  assign _3328_ = \u_csr.opcode_opcode_i [11:7] == 4'hd;
  assign _3329_ = \u_csr.opcode_opcode_i [11:7] == 4'hc;
  assign _3330_ = \u_csr.opcode_opcode_i [11:7] == 4'hb;
  assign _3331_ = \u_csr.opcode_opcode_i [11:7] == 4'ha;
  assign _3332_ = \u_csr.opcode_opcode_i [11:7] == 4'h9;
  assign _3333_ = \u_csr.opcode_opcode_i [11:7] == 4'h8;
  assign _3334_ = \u_csr.opcode_opcode_i [11:7] == 3'h7;
  assign _3335_ = \u_csr.opcode_opcode_i [11:7] == 3'h6;
  assign _3336_ = \u_csr.opcode_opcode_i [11:7] == 3'h5;
  assign _3337_ = \u_csr.opcode_opcode_i [11:7] == 3'h4;
  assign _3338_ = \u_csr.opcode_opcode_i [11:7] == 2'h3;
  assign _3339_ = \u_csr.opcode_opcode_i [11:7] == 2'h2;
  assign _3340_ = \u_csr.opcode_opcode_i [11:7] == 1'h1;
  assign _3341_ = ! \u_csr.opcode_opcode_i [11:7];
  logic [1:0] fangyuan200;
  assign fangyuan200 = { 1'h1, _3112_[29] };
  logic [1:0] fangyuan201;
  assign fangyuan201 = { _3312_, _3216_ };
  always @(1'hx or fangyuan200 or fangyuan201) begin
    casez (fangyuan201)
      2'b?1 :
        _3120_[29] = fangyuan200 [0:0] ;
      2'b1? :
        _3120_[29] = fangyuan200 [1:1] ;
      default:
        _3120_[29] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan202;
  assign fangyuan202 = { 1'h1, _3112_[27] };
  logic [1:0] fangyuan203;
  assign fangyuan203 = { _3314_, _3139_ };
  always @(1'hx or fangyuan202 or fangyuan203) begin
    casez (fangyuan203)
      2'b?1 :
        _3120_[27] = fangyuan202 [0:0] ;
      2'b1? :
        _3120_[27] = fangyuan202 [1:1] ;
      default:
        _3120_[27] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan204;
  assign fangyuan204 = { 1'h1, _3112_[25] };
  logic [1:0] fangyuan205;
  assign fangyuan205 = { _3316_, _3140_ };
  always @(1'hx or fangyuan204 or fangyuan205) begin
    casez (fangyuan205)
      2'b?1 :
        _3120_[25] = fangyuan204 [0:0] ;
      2'b1? :
        _3120_[25] = fangyuan204 [1:1] ;
      default:
        _3120_[25] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan206;
  assign fangyuan206 = { 1'h1, _3112_[23] };
  logic [1:0] fangyuan207;
  assign fangyuan207 = { _3318_, _3158_ };
  always @(1'hx or fangyuan206 or fangyuan207) begin
    casez (fangyuan207)
      2'b?1 :
        _3120_[23] = fangyuan206 [0:0] ;
      2'b1? :
        _3120_[23] = fangyuan206 [1:1] ;
      default:
        _3120_[23] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan208;
  assign fangyuan208 = { 1'h1, _3112_[21] };
  logic [1:0] fangyuan209;
  assign fangyuan209 = { _3320_, _3176_ };
  always @(1'hx or fangyuan208 or fangyuan209) begin
    casez (fangyuan209)
      2'b?1 :
        _3120_[21] = fangyuan208 [0:0] ;
      2'b1? :
        _3120_[21] = fangyuan208 [1:1] ;
      default:
        _3120_[21] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan210;
  assign fangyuan210 = { 1'h1, _3112_[19] };
  logic [1:0] fangyuan211;
  assign fangyuan211 = { _3322_, _3194_ };
  always @(1'hx or fangyuan210 or fangyuan211) begin
    casez (fangyuan211)
      2'b?1 :
        _3120_[19] = fangyuan210 [0:0] ;
      2'b1? :
        _3120_[19] = fangyuan210 [1:1] ;
      default:
        _3120_[19] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan212;
  assign fangyuan212 = { 1'h1, _3112_[17] };
  logic [1:0] fangyuan213;
  assign fangyuan213 = { _3324_, _3215_ };
  always @(1'hx or fangyuan212 or fangyuan213) begin
    casez (fangyuan213)
      2'b?1 :
        _3120_[17] = fangyuan212 [0:0] ;
      2'b1? :
        _3120_[17] = fangyuan212 [1:1] ;
      default:
        _3120_[17] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan214;
  assign fangyuan214 = { 1'h1, _3112_[15] };
  logic [1:0] fangyuan215;
  assign fangyuan215 = { _3326_, _3218_ };
  always @(1'hx or fangyuan214 or fangyuan215) begin
    casez (fangyuan215)
      2'b?1 :
        _3120_[15] = fangyuan214 [0:0] ;
      2'b1? :
        _3120_[15] = fangyuan214 [1:1] ;
      default:
        _3120_[15] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan216;
  assign fangyuan216 = { 1'h1, _3112_[13] };
  logic [1:0] fangyuan217;
  assign fangyuan217 = { _3328_, _3228_ };
  always @(1'hx or fangyuan216 or fangyuan217) begin
    casez (fangyuan217)
      2'b?1 :
        _3120_[13] = fangyuan216 [0:0] ;
      2'b1? :
        _3120_[13] = fangyuan216 [1:1] ;
      default:
        _3120_[13] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan218;
  assign fangyuan218 = { 1'h1, _3112_[11] };
  logic [1:0] fangyuan219;
  assign fangyuan219 = { _3330_, _3150_ };
  always @(1'hx or fangyuan218 or fangyuan219) begin
    casez (fangyuan219)
      2'b?1 :
        _3120_[11] = fangyuan218 [0:0] ;
      2'b1? :
        _3120_[11] = fangyuan218 [1:1] ;
      default:
        _3120_[11] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan220;
  assign fangyuan220 = { 1'h1, _3112_[9] };
  logic [1:0] fangyuan221;
  assign fangyuan221 = { _3332_, _3168_ };
  always @(1'hx or fangyuan220 or fangyuan221) begin
    casez (fangyuan221)
      2'b?1 :
        _3120_[9] = fangyuan220 [0:0] ;
      2'b1? :
        _3120_[9] = fangyuan220 [1:1] ;
      default:
        _3120_[9] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan222;
  assign fangyuan222 = { 1'h1, _3112_[7] };
  logic [1:0] fangyuan223;
  assign fangyuan223 = { _3334_, _3183_ };
  always @(1'hx or fangyuan222 or fangyuan223) begin
    casez (fangyuan223)
      2'b?1 :
        _3120_[7] = fangyuan222 [0:0] ;
      2'b1? :
        _3120_[7] = fangyuan222 [1:1] ;
      default:
        _3120_[7] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan224;
  assign fangyuan224 = { 1'h1, _3112_[5] };
  logic [1:0] fangyuan225;
  assign fangyuan225 = { _3336_, _3199_ };
  always @(1'hx or fangyuan224 or fangyuan225) begin
    casez (fangyuan225)
      2'b?1 :
        _3120_[5] = fangyuan224 [0:0] ;
      2'b1? :
        _3120_[5] = fangyuan224 [1:1] ;
      default:
        _3120_[5] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan226;
  assign fangyuan226 = { 1'h1, _3112_[3] };
  logic [1:0] fangyuan227;
  assign fangyuan227 = { _3338_, _3232_ };
  always @(1'hx or fangyuan226 or fangyuan227) begin
    casez (fangyuan227)
      2'b?1 :
        _3120_[3] = fangyuan226 [0:0] ;
      2'b1? :
        _3120_[3] = fangyuan226 [1:1] ;
      default:
        _3120_[3] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan228;
  assign fangyuan228 = { 1'h1, _3112_[1] };
  logic [1:0] fangyuan229;
  assign fangyuan229 = { _3340_, _3137_ };
  always @(1'hx or fangyuan228 or fangyuan229) begin
    casez (fangyuan229)
      2'b?1 :
        _3120_[1] = fangyuan228 [0:0] ;
      2'b1? :
        _3120_[1] = fangyuan228 [1:1] ;
      default:
        _3120_[1] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan230;
  assign fangyuan230 = { _3112_[31], 1'h1 };
  logic [1:0] fangyuan231;
  assign fangyuan231 = { _3227_, _3310_ };
  always @(1'hx or fangyuan230 or fangyuan231) begin
    casez (fangyuan231)
      2'b?1 :
        _3120_[31] = fangyuan230 [0:0] ;
      2'b1? :
        _3120_[31] = fangyuan230 [1:1] ;
      default:
        _3120_[31] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan232;
  assign fangyuan232 = { 1'h1, _3112_[26] };
  logic [1:0] fangyuan233;
  assign fangyuan233 = { _3315_, _3149_ };
  always @(1'hx or fangyuan232 or fangyuan233) begin
    casez (fangyuan233)
      2'b?1 :
        _3120_[26] = fangyuan232 [0:0] ;
      2'b1? :
        _3120_[26] = fangyuan232 [1:1] ;
      default:
        _3120_[26] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan234;
  assign fangyuan234 = { 1'h1, _3112_[22] };
  logic [1:0] fangyuan235;
  assign fangyuan235 = { _3319_, _3166_ };
  always @(1'hx or fangyuan234 or fangyuan235) begin
    casez (fangyuan235)
      2'b?1 :
        _3120_[22] = fangyuan234 [0:0] ;
      2'b1? :
        _3120_[22] = fangyuan234 [1:1] ;
      default:
        _3120_[22] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan236;
  assign fangyuan236 = { 1'h1, _3112_[18] };
  logic [1:0] fangyuan237;
  assign fangyuan237 = { _3323_, _3179_ };
  always @(1'hx or fangyuan236 or fangyuan237) begin
    casez (fangyuan237)
      2'b?1 :
        _3120_[18] = fangyuan236 [0:0] ;
      2'b1? :
        _3120_[18] = fangyuan236 [1:1] ;
      default:
        _3120_[18] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan238;
  assign fangyuan238 = { 1'h1, _3112_[14] };
  logic [1:0] fangyuan239;
  assign fangyuan239 = { _3327_, _3193_ };
  always @(1'hx or fangyuan238 or fangyuan239) begin
    casez (fangyuan239)
      2'b?1 :
        _3120_[14] = fangyuan238 [0:0] ;
      2'b1? :
        _3120_[14] = fangyuan238 [1:1] ;
      default:
        _3120_[14] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan240;
  assign fangyuan240 = { 1'h1, _3112_[10] };
  logic [1:0] fangyuan241;
  assign fangyuan241 = { _3331_, _3212_ };
  always @(1'hx or fangyuan240 or fangyuan241) begin
    casez (fangyuan241)
      2'b?1 :
        _3120_[10] = fangyuan240 [0:0] ;
      2'b1? :
        _3120_[10] = fangyuan240 [1:1] ;
      default:
        _3120_[10] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan242;
  assign fangyuan242 = { 1'h1, _3112_[6] };
  logic [1:0] fangyuan243;
  assign fangyuan243 = { _3335_, _3230_ };
  always @(1'hx or fangyuan242 or fangyuan243) begin
    casez (fangyuan243)
      2'b?1 :
        _3120_[6] = fangyuan242 [0:0] ;
      2'b1? :
        _3120_[6] = fangyuan242 [1:1] ;
      default:
        _3120_[6] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan244;
  assign fangyuan244 = { 1'h1, _3112_[2] };
  logic [1:0] fangyuan245;
  assign fangyuan245 = { _3339_, _3146_ };
  always @(1'hx or fangyuan244 or fangyuan245) begin
    casez (fangyuan245)
      2'b?1 :
        _3120_[2] = fangyuan244 [0:0] ;
      2'b1? :
        _3120_[2] = fangyuan244 [1:1] ;
      default:
        _3120_[2] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan246;
  assign fangyuan246 = { 1'h1, _3112_[28] };
  logic [1:0] fangyuan247;
  assign fangyuan247 = { _3313_, _3231_ };
  always @(1'hx or fangyuan246 or fangyuan247) begin
    casez (fangyuan247)
      2'b?1 :
        _3120_[28] = fangyuan246 [0:0] ;
      2'b1? :
        _3120_[28] = fangyuan246 [1:1] ;
      default:
        _3120_[28] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan248;
  assign fangyuan248 = { 1'h1, _3112_[20] };
  logic [1:0] fangyuan249;
  assign fangyuan249 = { _3321_, _3148_ };
  always @(1'hx or fangyuan248 or fangyuan249) begin
    casez (fangyuan249)
      2'b?1 :
        _3120_[20] = fangyuan248 [0:0] ;
      2'b1? :
        _3120_[20] = fangyuan248 [1:1] ;
      default:
        _3120_[20] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan250;
  assign fangyuan250 = { 1'h1, _3112_[12] };
  logic [1:0] fangyuan251;
  assign fangyuan251 = { _3329_, _3160_ };
  always @(1'hx or fangyuan250 or fangyuan251) begin
    casez (fangyuan251)
      2'b?1 :
        _3120_[12] = fangyuan250 [0:0] ;
      2'b1? :
        _3120_[12] = fangyuan250 [1:1] ;
      default:
        _3120_[12] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan252;
  assign fangyuan252 = { 1'h1, _3112_[4] };
  logic [1:0] fangyuan253;
  assign fangyuan253 = { _3337_, _3177_ };
  always @(1'hx or fangyuan252 or fangyuan253) begin
    casez (fangyuan253)
      2'b?1 :
        _3120_[4] = fangyuan252 [0:0] ;
      2'b1? :
        _3120_[4] = fangyuan252 [1:1] ;
      default:
        _3120_[4] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan254;
  assign fangyuan254 = { 1'h1, _3112_[24] };
  logic [1:0] fangyuan255;
  assign fangyuan255 = { _3317_, _3187_ };
  always @(1'hx or fangyuan254 or fangyuan255) begin
    casez (fangyuan255)
      2'b?1 :
        _3120_[24] = fangyuan254 [0:0] ;
      2'b1? :
        _3120_[24] = fangyuan254 [1:1] ;
      default:
        _3120_[24] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan256;
  assign fangyuan256 = { 1'h1, _3112_[8] };
  logic [1:0] fangyuan257;
  assign fangyuan257 = { _3333_, _3203_ };
  always @(1'hx or fangyuan256 or fangyuan257) begin
    casez (fangyuan257)
      2'b?1 :
        _3120_[8] = fangyuan256 [0:0] ;
      2'b1? :
        _3120_[8] = fangyuan256 [1:1] ;
      default:
        _3120_[8] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan258;
  assign fangyuan258 = { 1'h1, _3112_[16] };
  logic [1:0] fangyuan259;
  assign fangyuan259 = { _3325_, _3220_ };
  always @(1'hx or fangyuan258 or fangyuan259) begin
    casez (fangyuan259)
      2'b?1 :
        _3120_[16] = fangyuan258 [0:0] ;
      2'b1? :
        _3120_[16] = fangyuan258 [1:1] ;
      default:
        _3120_[16] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan260;
  assign fangyuan260 = { 1'h1, _3112_[0] };
  logic [1:0] fangyuan261;
  assign fangyuan261 = { _3341_, _3172_ };
  always @(1'hx or fangyuan260 or fangyuan261) begin
    casez (fangyuan261)
      2'b?1 :
        _3120_[0] = fangyuan260 [0:0] ;
      2'b1? :
        _3120_[0] = fangyuan260 [1:1] ;
      default:
        _3120_[0] = 1'hx ;
    endcase
  end
  assign _3119_ = _3276_ ? _3120_ : _3112_;
  assign _3118_ = _3275_ ? _3119_ : _3112_;
  assign _3084_ = _3275_ ? 1'h1 : 1'h0;
  assign _3117_ = _3296_ ? _3112_ : _3118_;
  assign \u_div.opcode_valid_i = _3296_ ? 1'h0 : _3084_;
  assign _3112_ = _3274_ ? 32'hffffffff : _3100_;
  logic [1:0] fangyuan262;
  assign fangyuan262 = { 1'h1, _3078_[30] };
  logic [1:0] fangyuan263;
  assign fangyuan263 = { _3343_, _3175_ };
  always @(1'hx or fangyuan262 or fangyuan263) begin
    casez (fangyuan263)
      2'b?1 :
        _3107_[30] = fangyuan262 [0:0] ;
      2'b1? :
        _3107_[30] = fangyuan262 [1:1] ;
      default:
        _3107_[30] = 1'hx ;
    endcase
  end
  assign _3342_ = \u_issue.pipe1_rd_e1_w == 5'h1f;
  assign _3343_ = \u_issue.pipe1_rd_e1_w == 5'h1e;
  assign _3344_ = \u_issue.pipe1_rd_e1_w == 5'h1d;
  assign _3345_ = \u_issue.pipe1_rd_e1_w == 5'h1c;
  assign _3346_ = \u_issue.pipe1_rd_e1_w == 5'h1b;
  assign _3347_ = \u_issue.pipe1_rd_e1_w == 5'h1a;
  assign _3348_ = \u_issue.pipe1_rd_e1_w == 5'h19;
  assign _3349_ = \u_issue.pipe1_rd_e1_w == 5'h18;
  assign _3350_ = \u_issue.pipe1_rd_e1_w == 5'h17;
  assign _3351_ = \u_issue.pipe1_rd_e1_w == 5'h16;
  assign _3352_ = \u_issue.pipe1_rd_e1_w == 5'h15;
  assign _3353_ = \u_issue.pipe1_rd_e1_w == 5'h14;
  assign _3354_ = \u_issue.pipe1_rd_e1_w == 5'h13;
  assign _3355_ = \u_issue.pipe1_rd_e1_w == 5'h12;
  assign _3356_ = \u_issue.pipe1_rd_e1_w == 5'h11;
  assign _3357_ = \u_issue.pipe1_rd_e1_w == 5'h10;
  assign _3358_ = \u_issue.pipe1_rd_e1_w == 4'hf;
  assign _3359_ = \u_issue.pipe1_rd_e1_w == 4'he;
  assign _3360_ = \u_issue.pipe1_rd_e1_w == 4'hd;
  assign _3361_ = \u_issue.pipe1_rd_e1_w == 4'hc;
  assign _3362_ = \u_issue.pipe1_rd_e1_w == 4'hb;
  assign _3363_ = \u_issue.pipe1_rd_e1_w == 4'ha;
  assign _3364_ = \u_issue.pipe1_rd_e1_w == 4'h9;
  assign _3365_ = \u_issue.pipe1_rd_e1_w == 4'h8;
  assign _3366_ = \u_issue.pipe1_rd_e1_w == 3'h7;
  assign _3367_ = \u_issue.pipe1_rd_e1_w == 3'h6;
  assign _3368_ = \u_issue.pipe1_rd_e1_w == 3'h5;
  assign _3369_ = \u_issue.pipe1_rd_e1_w == 3'h4;
  assign _3370_ = \u_issue.pipe1_rd_e1_w == 2'h3;
  assign _3371_ = \u_issue.pipe1_rd_e1_w == 2'h2;
  assign _3372_ = \u_issue.pipe1_rd_e1_w == 1'h1;
  assign _3373_ = ! \u_issue.pipe1_rd_e1_w ;
  logic [1:0] fangyuan264;
  assign fangyuan264 = { 1'h1, _3078_[29] };
  logic [1:0] fangyuan265;
  assign fangyuan265 = { _3344_, _3204_ };
  always @(1'hx or fangyuan264 or fangyuan265) begin
    casez (fangyuan265)
      2'b?1 :
        _3107_[29] = fangyuan264 [0:0] ;
      2'b1? :
        _3107_[29] = fangyuan264 [1:1] ;
      default:
        _3107_[29] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan266;
  assign fangyuan266 = { 1'h1, _3078_[27] };
  logic [1:0] fangyuan267;
  assign fangyuan267 = { _3346_, _3138_ };
  always @(1'hx or fangyuan266 or fangyuan267) begin
    casez (fangyuan267)
      2'b?1 :
        _3107_[27] = fangyuan266 [0:0] ;
      2'b1? :
        _3107_[27] = fangyuan266 [1:1] ;
      default:
        _3107_[27] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan268;
  assign fangyuan268 = { 1'h1, _3078_[25] };
  logic [1:0] fangyuan269;
  assign fangyuan269 = { _3348_, _3147_ };
  always @(1'hx or fangyuan268 or fangyuan269) begin
    casez (fangyuan269)
      2'b?1 :
        _3107_[25] = fangyuan268 [0:0] ;
      2'b1? :
        _3107_[25] = fangyuan268 [1:1] ;
      default:
        _3107_[25] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan270;
  assign fangyuan270 = { 1'h1, _3078_[23] };
  logic [1:0] fangyuan271;
  assign fangyuan271 = { _3350_, _3159_ };
  always @(1'hx or fangyuan270 or fangyuan271) begin
    casez (fangyuan271)
      2'b?1 :
        _3107_[23] = fangyuan270 [0:0] ;
      2'b1? :
        _3107_[23] = fangyuan270 [1:1] ;
      default:
        _3107_[23] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan272;
  assign fangyuan272 = { 1'h1, _3078_[21] };
  logic [1:0] fangyuan273;
  assign fangyuan273 = { _3352_, _3169_ };
  always @(1'hx or fangyuan272 or fangyuan273) begin
    casez (fangyuan273)
      2'b?1 :
        _3107_[21] = fangyuan272 [0:0] ;
      2'b1? :
        _3107_[21] = fangyuan272 [1:1] ;
      default:
        _3107_[21] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan274;
  assign fangyuan274 = { 1'h1, _3078_[19] };
  logic [1:0] fangyuan275;
  assign fangyuan275 = { _3354_, _3185_ };
  always @(1'hx or fangyuan274 or fangyuan275) begin
    casez (fangyuan275)
      2'b?1 :
        _3107_[19] = fangyuan274 [0:0] ;
      2'b1? :
        _3107_[19] = fangyuan274 [1:1] ;
      default:
        _3107_[19] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan276;
  assign fangyuan276 = { 1'h1, _3078_[17] };
  logic [1:0] fangyuan277;
  assign fangyuan277 = { _3356_, _3196_ };
  always @(1'hx or fangyuan276 or fangyuan277) begin
    casez (fangyuan277)
      2'b?1 :
        _3107_[17] = fangyuan276 [0:0] ;
      2'b1? :
        _3107_[17] = fangyuan276 [1:1] ;
      default:
        _3107_[17] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan278;
  assign fangyuan278 = { 1'h1, _3078_[15] };
  logic [1:0] fangyuan279;
  assign fangyuan279 = { _3358_, _3210_ };
  always @(1'hx or fangyuan278 or fangyuan279) begin
    casez (fangyuan279)
      2'b?1 :
        _3107_[15] = fangyuan278 [0:0] ;
      2'b1? :
        _3107_[15] = fangyuan278 [1:1] ;
      default:
        _3107_[15] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan280;
  assign fangyuan280 = { 1'h1, _3078_[13] };
  logic [1:0] fangyuan281;
  assign fangyuan281 = { _3360_, _3156_ };
  always @(1'hx or fangyuan280 or fangyuan281) begin
    casez (fangyuan281)
      2'b?1 :
        _3107_[13] = fangyuan280 [0:0] ;
      2'b1? :
        _3107_[13] = fangyuan280 [1:1] ;
      default:
        _3107_[13] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan282;
  assign fangyuan282 = { 1'h1, _3078_[11] };
  logic [1:0] fangyuan283;
  assign fangyuan283 = { _3362_, _3223_ };
  always @(1'hx or fangyuan282 or fangyuan283) begin
    casez (fangyuan283)
      2'b?1 :
        _3107_[11] = fangyuan282 [0:0] ;
      2'b1? :
        _3107_[11] = fangyuan282 [1:1] ;
      default:
        _3107_[11] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan284;
  assign fangyuan284 = { 1'h1, _3078_[9] };
  logic [1:0] fangyuan285;
  assign fangyuan285 = { _3364_, _3162_ };
  always @(1'hx or fangyuan284 or fangyuan285) begin
    casez (fangyuan285)
      2'b?1 :
        _3107_[9] = fangyuan284 [0:0] ;
      2'b1? :
        _3107_[9] = fangyuan284 [1:1] ;
      default:
        _3107_[9] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan286;
  assign fangyuan286 = { 1'h1, _3078_[7] };
  logic [1:0] fangyuan287;
  assign fangyuan287 = { _3366_, _3192_ };
  always @(1'hx or fangyuan286 or fangyuan287) begin
    casez (fangyuan287)
      2'b?1 :
        _3107_[7] = fangyuan286 [0:0] ;
      2'b1? :
        _3107_[7] = fangyuan286 [1:1] ;
      default:
        _3107_[7] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan288;
  assign fangyuan288 = { 1'h1, _3078_[5] };
  logic [1:0] fangyuan289;
  assign fangyuan289 = { _3368_, _3224_ };
  always @(1'hx or fangyuan288 or fangyuan289) begin
    casez (fangyuan289)
      2'b?1 :
        _3107_[5] = fangyuan288 [0:0] ;
      2'b1? :
        _3107_[5] = fangyuan288 [1:1] ;
      default:
        _3107_[5] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan290;
  assign fangyuan290 = { 1'h1, _3078_[3] };
  logic [1:0] fangyuan291;
  assign fangyuan291 = { _3370_, _3143_ };
  always @(1'hx or fangyuan290 or fangyuan291) begin
    casez (fangyuan291)
      2'b?1 :
        _3107_[3] = fangyuan290 [0:0] ;
      2'b1? :
        _3107_[3] = fangyuan290 [1:1] ;
      default:
        _3107_[3] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan292;
  assign fangyuan292 = { 1'h1, _3078_[1] };
  logic [1:0] fangyuan293;
  assign fangyuan293 = { _3372_, _3154_ };
  always @(1'hx or fangyuan292 or fangyuan293) begin
    casez (fangyuan293)
      2'b?1 :
        _3107_[1] = fangyuan292 [0:0] ;
      2'b1? :
        _3107_[1] = fangyuan292 [1:1] ;
      default:
        _3107_[1] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan294;
  assign fangyuan294 = { _3078_[31], 1'h1 };
  logic [1:0] fangyuan295;
  assign fangyuan295 = { _3167_, _3342_ };
  always @(1'hx or fangyuan294 or fangyuan295) begin
    casez (fangyuan295)
      2'b?1 :
        _3107_[31] = fangyuan294 [0:0] ;
      2'b1? :
        _3107_[31] = fangyuan294 [1:1] ;
      default:
        _3107_[31] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan296;
  assign fangyuan296 = { 1'h1, _3078_[26] };
  logic [1:0] fangyuan297;
  assign fangyuan297 = { _3347_, _3178_ };
  always @(1'hx or fangyuan296 or fangyuan297) begin
    casez (fangyuan297)
      2'b?1 :
        _3107_[26] = fangyuan296 [0:0] ;
      2'b1? :
        _3107_[26] = fangyuan296 [1:1] ;
      default:
        _3107_[26] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan298;
  assign fangyuan298 = { 1'h1, _3078_[22] };
  logic [1:0] fangyuan299;
  assign fangyuan299 = { _3351_, _3186_ };
  always @(1'hx or fangyuan298 or fangyuan299) begin
    casez (fangyuan299)
      2'b?1 :
        _3107_[22] = fangyuan298 [0:0] ;
      2'b1? :
        _3107_[22] = fangyuan298 [1:1] ;
      default:
        _3107_[22] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan300;
  assign fangyuan300 = { 1'h1, _3078_[18] };
  logic [1:0] fangyuan301;
  assign fangyuan301 = { _3355_, _3198_ };
  always @(1'hx or fangyuan300 or fangyuan301) begin
    casez (fangyuan301)
      2'b?1 :
        _3107_[18] = fangyuan300 [0:0] ;
      2'b1? :
        _3107_[18] = fangyuan300 [1:1] ;
      default:
        _3107_[18] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan302;
  assign fangyuan302 = { 1'h1, _3078_[14] };
  logic [1:0] fangyuan303;
  assign fangyuan303 = { _3359_, _3213_ };
  always @(1'hx or fangyuan302 or fangyuan303) begin
    casez (fangyuan303)
      2'b?1 :
        _3107_[14] = fangyuan302 [0:0] ;
      2'b1? :
        _3107_[14] = fangyuan302 [1:1] ;
      default:
        _3107_[14] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan304;
  assign fangyuan304 = { 1'h1, _3078_[10] };
  logic [1:0] fangyuan305;
  assign fangyuan305 = { _3363_, _3221_ };
  always @(1'hx or fangyuan304 or fangyuan305) begin
    casez (fangyuan305)
      2'b?1 :
        _3107_[10] = fangyuan304 [0:0] ;
      2'b1? :
        _3107_[10] = fangyuan304 [1:1] ;
      default:
        _3107_[10] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan306;
  assign fangyuan306 = { 1'h1, _3078_[6] };
  logic [1:0] fangyuan307;
  assign fangyuan307 = { _3367_, _3226_ };
  always @(1'hx or fangyuan306 or fangyuan307) begin
    casez (fangyuan307)
      2'b?1 :
        _3107_[6] = fangyuan306 [0:0] ;
      2'b1? :
        _3107_[6] = fangyuan306 [1:1] ;
      default:
        _3107_[6] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan308;
  assign fangyuan308 = { 1'h1, _3078_[2] };
  logic [1:0] fangyuan309;
  assign fangyuan309 = { _3371_, _3165_ };
  always @(1'hx or fangyuan308 or fangyuan309) begin
    casez (fangyuan309)
      2'b?1 :
        _3107_[2] = fangyuan308 [0:0] ;
      2'b1? :
        _3107_[2] = fangyuan308 [1:1] ;
      default:
        _3107_[2] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan310;
  assign fangyuan310 = { 1'h1, _3078_[28] };
  logic [1:0] fangyuan311;
  assign fangyuan311 = { _3345_, _3190_ };
  always @(1'hx or fangyuan310 or fangyuan311) begin
    casez (fangyuan311)
      2'b?1 :
        _3107_[28] = fangyuan310 [0:0] ;
      2'b1? :
        _3107_[28] = fangyuan310 [1:1] ;
      default:
        _3107_[28] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan312;
  assign fangyuan312 = { 1'h1, _3078_[20] };
  logic [1:0] fangyuan313;
  assign fangyuan313 = { _3353_, _3222_ };
  always @(1'hx or fangyuan312 or fangyuan313) begin
    casez (fangyuan313)
      2'b?1 :
        _3107_[20] = fangyuan312 [0:0] ;
      2'b1? :
        _3107_[20] = fangyuan312 [1:1] ;
      default:
        _3107_[20] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan314;
  assign fangyuan314 = { 1'h1, _3078_[12] };
  logic [1:0] fangyuan315;
  assign fangyuan315 = { _3361_, _3141_ };
  always @(1'hx or fangyuan314 or fangyuan315) begin
    casez (fangyuan315)
      2'b?1 :
        _3107_[12] = fangyuan314 [0:0] ;
      2'b1? :
        _3107_[12] = fangyuan314 [1:1] ;
      default:
        _3107_[12] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan316;
  assign fangyuan316 = { 1'h1, _3078_[4] };
  logic [1:0] fangyuan317;
  assign fangyuan317 = { _3369_, _3151_ };
  always @(1'hx or fangyuan316 or fangyuan317) begin
    casez (fangyuan317)
      2'b?1 :
        _3107_[4] = fangyuan316 [0:0] ;
      2'b1? :
        _3107_[4] = fangyuan316 [1:1] ;
      default:
        _3107_[4] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan318;
  assign fangyuan318 = { 1'h1, _3078_[24] };
  logic [1:0] fangyuan319;
  assign fangyuan319 = { _3349_, _3164_ };
  always @(1'hx or fangyuan318 or fangyuan319) begin
    casez (fangyuan319)
      2'b?1 :
        _3107_[24] = fangyuan318 [0:0] ;
      2'b1? :
        _3107_[24] = fangyuan318 [1:1] ;
      default:
        _3107_[24] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan320;
  assign fangyuan320 = { 1'h1, _3078_[8] };
  logic [1:0] fangyuan321;
  assign fangyuan321 = { _3365_, _3174_ };
  always @(1'hx or fangyuan320 or fangyuan321) begin
    casez (fangyuan321)
      2'b?1 :
        _3107_[8] = fangyuan320 [0:0] ;
      2'b1? :
        _3107_[8] = fangyuan320 [1:1] ;
      default:
        _3107_[8] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan322;
  assign fangyuan322 = { 1'h1, _3078_[16] };
  logic [1:0] fangyuan323;
  assign fangyuan323 = { _3357_, _3184_ };
  always @(1'hx or fangyuan322 or fangyuan323) begin
    casez (fangyuan323)
      2'b?1 :
        _3107_[16] = fangyuan322 [0:0] ;
      2'b1? :
        _3107_[16] = fangyuan322 [1:1] ;
      default:
        _3107_[16] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan324;
  assign fangyuan324 = { 1'h1, _3078_[0] };
  logic [1:0] fangyuan325;
  assign fangyuan325 = { _3373_, _3195_ };
  always @(1'hx or fangyuan324 or fangyuan325) begin
    casez (fangyuan325)
      2'b?1 :
        _3107_[0] = fangyuan324 [0:0] ;
      2'b1? :
        _3107_[0] = fangyuan324 [1:1] ;
      default:
        _3107_[0] = 1'hx ;
    endcase
  end
  assign _3100_ = _3288_ ? _3107_ : _3078_;
  logic [1:0] fangyuan326;
  assign fangyuan326 = { _3375_, _3205_ };
  always @(1'hx or fangyuan326) begin
    casez (fangyuan326)
      2'b?1 :
        _3092_[30] = 1'b0 ;
      2'b1? :
        _3092_[30] = 1'b1 ;
      default:
        _3092_[30] = 1'hx ;
    endcase
  end
  assign _3374_ = \u_issue.pipe0_rd_e1_w == 5'h1f;
  assign _3375_ = \u_issue.pipe0_rd_e1_w == 5'h1e;
  assign _3376_ = \u_issue.pipe0_rd_e1_w == 5'h1d;
  assign _3377_ = \u_issue.pipe0_rd_e1_w == 5'h1c;
  assign _3378_ = \u_issue.pipe0_rd_e1_w == 5'h1b;
  assign _3379_ = \u_issue.pipe0_rd_e1_w == 5'h1a;
  assign _3380_ = \u_issue.pipe0_rd_e1_w == 5'h19;
  assign _3381_ = \u_issue.pipe0_rd_e1_w == 5'h18;
  assign _3382_ = \u_issue.pipe0_rd_e1_w == 5'h17;
  assign _3383_ = \u_issue.pipe0_rd_e1_w == 5'h16;
  assign _3384_ = \u_issue.pipe0_rd_e1_w == 5'h15;
  assign _3385_ = \u_issue.pipe0_rd_e1_w == 5'h14;
  assign _3386_ = \u_issue.pipe0_rd_e1_w == 5'h13;
  assign _3387_ = \u_issue.pipe0_rd_e1_w == 5'h12;
  assign _3388_ = \u_issue.pipe0_rd_e1_w == 5'h11;
  assign _3389_ = \u_issue.pipe0_rd_e1_w == 5'h10;
  assign _3390_ = \u_issue.pipe0_rd_e1_w == 4'hf;
  assign _3391_ = \u_issue.pipe0_rd_e1_w == 4'he;
  assign _3392_ = \u_issue.pipe0_rd_e1_w == 4'hd;
  assign _3393_ = \u_issue.pipe0_rd_e1_w == 4'hc;
  assign _3394_ = \u_issue.pipe0_rd_e1_w == 4'hb;
  assign _3395_ = \u_issue.pipe0_rd_e1_w == 4'ha;
  assign _3396_ = \u_issue.pipe0_rd_e1_w == 4'h9;
  assign _3397_ = \u_issue.pipe0_rd_e1_w == 4'h8;
  assign _3398_ = \u_issue.pipe0_rd_e1_w == 3'h7;
  assign _3399_ = \u_issue.pipe0_rd_e1_w == 3'h6;
  assign _3400_ = \u_issue.pipe0_rd_e1_w == 3'h5;
  assign _3401_ = \u_issue.pipe0_rd_e1_w == 3'h4;
  assign _3402_ = \u_issue.pipe0_rd_e1_w == 2'h3;
  assign _3403_ = \u_issue.pipe0_rd_e1_w == 2'h2;
  assign _3404_ = \u_issue.pipe0_rd_e1_w == 1'h1;
  assign _3405_ = ! \u_issue.pipe0_rd_e1_w ;
  logic [1:0] fangyuan327;
  assign fangyuan327 = { _3376_, _3209_ };
  always @(1'hx or fangyuan327) begin
    casez (fangyuan327)
      2'b?1 :
        _3092_[29] = 1'b0 ;
      2'b1? :
        _3092_[29] = 1'b1 ;
      default:
        _3092_[29] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan328;
  assign fangyuan328 = { _3378_, _3219_ };
  always @(1'hx or fangyuan328) begin
    casez (fangyuan328)
      2'b?1 :
        _3092_[27] = 1'b0 ;
      2'b1? :
        _3092_[27] = 1'b1 ;
      default:
        _3092_[27] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan329;
  assign fangyuan329 = { _3380_, _3157_ };
  always @(1'hx or fangyuan329) begin
    casez (fangyuan329)
      2'b?1 :
        _3092_[25] = 1'b0 ;
      2'b1? :
        _3092_[25] = 1'b1 ;
      default:
        _3092_[25] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan330;
  assign fangyuan330 = { _3382_, _3144_ };
  always @(1'hx or fangyuan330) begin
    casez (fangyuan330)
      2'b?1 :
        _3092_[23] = 1'b0 ;
      2'b1? :
        _3092_[23] = 1'b1 ;
      default:
        _3092_[23] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan331;
  assign fangyuan331 = { _3384_, _3173_ };
  always @(1'hx or fangyuan331) begin
    casez (fangyuan331)
      2'b?1 :
        _3092_[21] = 1'b0 ;
      2'b1? :
        _3092_[21] = 1'b1 ;
      default:
        _3092_[21] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan332;
  assign fangyuan332 = { _3386_, _3197_ };
  always @(1'hx or fangyuan332) begin
    casez (fangyuan332)
      2'b?1 :
        _3092_[19] = 1'b0 ;
      2'b1? :
        _3092_[19] = 1'b1 ;
      default:
        _3092_[19] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan333;
  assign fangyuan333 = { _3388_, _3225_ };
  always @(1'hx or fangyuan333) begin
    casez (fangyuan333)
      2'b?1 :
        _3092_[17] = 1'b0 ;
      2'b1? :
        _3092_[17] = 1'b1 ;
      default:
        _3092_[17] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan334;
  assign fangyuan334 = { _3390_, _3142_ };
  always @(1'hx or fangyuan334) begin
    casez (fangyuan334)
      2'b?1 :
        _3092_[15] = 1'b0 ;
      2'b1? :
        _3092_[15] = 1'b1 ;
      default:
        _3092_[15] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan335;
  assign fangyuan335 = { _3392_, _3152_ };
  always @(1'hx or fangyuan335) begin
    casez (fangyuan335)
      2'b?1 :
        _3092_[13] = 1'b0 ;
      2'b1? :
        _3092_[13] = 1'b1 ;
      default:
        _3092_[13] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan336;
  assign fangyuan336 = { _3394_, _3161_ };
  always @(1'hx or fangyuan336) begin
    casez (fangyuan336)
      2'b?1 :
        _3092_[11] = 1'b0 ;
      2'b1? :
        _3092_[11] = 1'b1 ;
      default:
        _3092_[11] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan337;
  assign fangyuan337 = { _3396_, _3171_ };
  always @(1'hx or fangyuan337) begin
    casez (fangyuan337)
      2'b?1 :
        _3092_[9] = 1'b0 ;
      2'b1? :
        _3092_[9] = 1'b1 ;
      default:
        _3092_[9] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan338;
  assign fangyuan338 = { _3398_, _3181_ };
  always @(1'hx or fangyuan338) begin
    casez (fangyuan338)
      2'b?1 :
        _3092_[7] = 1'b0 ;
      2'b1? :
        _3092_[7] = 1'b1 ;
      default:
        _3092_[7] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan339;
  assign fangyuan339 = { _3400_, _3191_ };
  always @(1'hx or fangyuan339) begin
    casez (fangyuan339)
      2'b?1 :
        _3092_[5] = 1'b0 ;
      2'b1? :
        _3092_[5] = 1'b1 ;
      default:
        _3092_[5] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan340;
  assign fangyuan340 = { _3402_, _3202_ };
  always @(1'hx or fangyuan340) begin
    casez (fangyuan340)
      2'b?1 :
        _3092_[3] = 1'b0 ;
      2'b1? :
        _3092_[3] = 1'b1 ;
      default:
        _3092_[3] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan341;
  assign fangyuan341 = { _3404_, _3207_ };
  always @(1'hx or fangyuan341) begin
    casez (fangyuan341)
      2'b?1 :
        _3092_[1] = 1'b0 ;
      2'b1? :
        _3092_[1] = 1'b1 ;
      default:
        _3092_[1] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan342;
  assign fangyuan342 = { _3214_, _3374_ };
  always @(1'hx or fangyuan342) begin
    casez (fangyuan342)
      2'b?1 :
        _3092_[31] = 1'b1 ;
      2'b1? :
        _3092_[31] = 1'b0 ;
      default:
        _3092_[31] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan343;
  assign fangyuan343 = { _3379_, _3201_ };
  always @(1'hx or fangyuan343) begin
    casez (fangyuan343)
      2'b?1 :
        _3092_[26] = 1'b0 ;
      2'b1? :
        _3092_[26] = 1'b1 ;
      default:
        _3092_[26] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan344;
  assign fangyuan344 = { _3383_, _3217_ };
  always @(1'hx or fangyuan344) begin
    casez (fangyuan344)
      2'b?1 :
        _3092_[22] = 1'b0 ;
      2'b1? :
        _3092_[22] = 1'b1 ;
      default:
        _3092_[22] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan345;
  assign fangyuan345 = { _3387_, _3155_ };
  always @(1'hx or fangyuan345) begin
    casez (fangyuan345)
      2'b?1 :
        _3092_[18] = 1'b0 ;
      2'b1? :
        _3092_[18] = 1'b1 ;
      default:
        _3092_[18] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan346;
  assign fangyuan346 = { _3391_, _3182_ };
  always @(1'hx or fangyuan346) begin
    casez (fangyuan346)
      2'b?1 :
        _3092_[14] = 1'b0 ;
      2'b1? :
        _3092_[14] = 1'b1 ;
      default:
        _3092_[14] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan347;
  assign fangyuan347 = { _3395_, _3208_ };
  always @(1'hx or fangyuan347) begin
    casez (fangyuan347)
      2'b?1 :
        _3092_[10] = 1'b0 ;
      2'b1? :
        _3092_[10] = 1'b1 ;
      default:
        _3092_[10] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan348;
  assign fangyuan348 = { _3399_, _3229_ };
  always @(1'hx or fangyuan348) begin
    casez (fangyuan348)
      2'b?1 :
        _3092_[6] = 1'b0 ;
      2'b1? :
        _3092_[6] = 1'b1 ;
      default:
        _3092_[6] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan349;
  assign fangyuan349 = { _3403_, _3145_ };
  always @(1'hx or fangyuan349) begin
    casez (fangyuan349)
      2'b?1 :
        _3092_[2] = 1'b0 ;
      2'b1? :
        _3092_[2] = 1'b1 ;
      default:
        _3092_[2] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan350;
  assign fangyuan350 = { _3377_, _3153_ };
  always @(1'hx or fangyuan350) begin
    casez (fangyuan350)
      2'b?1 :
        _3092_[28] = 1'b0 ;
      2'b1? :
        _3092_[28] = 1'b1 ;
      default:
        _3092_[28] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan351;
  assign fangyuan351 = { _3385_, _3163_ };
  always @(1'hx or fangyuan351) begin
    casez (fangyuan351)
      2'b?1 :
        _3092_[20] = 1'b0 ;
      2'b1? :
        _3092_[20] = 1'b1 ;
      default:
        _3092_[20] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan352;
  assign fangyuan352 = { _3393_, _3170_ };
  always @(1'hx or fangyuan352) begin
    casez (fangyuan352)
      2'b?1 :
        _3092_[12] = 1'b0 ;
      2'b1? :
        _3092_[12] = 1'b1 ;
      default:
        _3092_[12] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan353;
  assign fangyuan353 = { _3401_, _3180_ };
  always @(1'hx or fangyuan353) begin
    casez (fangyuan353)
      2'b?1 :
        _3092_[4] = 1'b0 ;
      2'b1? :
        _3092_[4] = 1'b1 ;
      default:
        _3092_[4] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan354;
  assign fangyuan354 = { _3381_, _3189_ };
  always @(1'hx or fangyuan354) begin
    casez (fangyuan354)
      2'b?1 :
        _3092_[24] = 1'b0 ;
      2'b1? :
        _3092_[24] = 1'b1 ;
      default:
        _3092_[24] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan355;
  assign fangyuan355 = { _3397_, _3200_ };
  always @(1'hx or fangyuan355) begin
    casez (fangyuan355)
      2'b?1 :
        _3092_[8] = 1'b0 ;
      2'b1? :
        _3092_[8] = 1'b1 ;
      default:
        _3092_[8] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan356;
  assign fangyuan356 = { _3389_, _3206_ };
  always @(1'hx or fangyuan356) begin
    casez (fangyuan356)
      2'b?1 :
        _3092_[16] = 1'b0 ;
      2'b1? :
        _3092_[16] = 1'b1 ;
      default:
        _3092_[16] = 1'hx ;
    endcase
  end
  logic [1:0] fangyuan357;
  assign fangyuan357 = { _3405_, _3211_ };
  always @(1'hx or fangyuan357) begin
    casez (fangyuan357)
      2'b?1 :
        _3092_[0] = 1'b0 ;
      2'b1? :
        _3092_[0] = 1'b1 ;
      default:
        _3092_[0] = 1'hx ;
    endcase
  end
  assign _3078_ = _3287_ ? _3092_ : 32'h00000000;
  assign _3406_ = \u_issue.pipe0_csr_wb_w ? 1'h0 : \u_issue.csr_pending_q ;
  assign _3407_ = _3268_ ? 1'h1 : _3406_;
  assign _3408_ = \u_issue.squash_w ? 1'h0 : _3407_;
  assign _3071_ = rst_i ? 1'h0 : _3408_;
  assign _3409_ = \u_div.valid_q ? 1'h0 : \u_issue.div_pending_q ;
  assign _3410_ = _3267_ ? 1'h1 : _3409_;
  assign _3411_ = \u_issue.squash_w ? 1'h0 : _3410_;
  assign _3072_ = rst_i ? 1'h0 : _3411_;
  assign _3085_ = \u_issue.slot1_valid_r ? \u_frontend.u_decode.u_fifo.info1_out_o : 2'h0;
  logic [31:0] fangyuan358;
  assign fangyuan358 = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign _3086_ = \u_issue.slot1_valid_r ? fangyuan358 : 32'h00000000;
  assign _3087_ = \u_issue.slot1_valid_r ? \u_frontend.u_decode.u_fifo.data1_out_o : 32'h00000000;
  assign _3088_ = \u_issue.slot1_valid_r ? 1'h1 : 1'h0;
  assign \u_issue.opcode_b_fault_r = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_fifo.info1_out_o : 2'h0;
  logic [31:0] fangyuan359;
  assign fangyuan359 = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign \u_exec1.opcode_pc_i = \u_issue.slot0_valid_r ? fangyuan359 : 32'h00000000;
  assign \u_exec1.opcode_opcode_i = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_fifo.data1_out_o : 32'h00000000;
  assign \u_issue.opcode_a_fault_r = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_fifo.info0_out_o : _3085_;
  logic [31:0] fangyuan360;
  assign fangyuan360 = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h0 };
  assign \u_exec0.opcode_pc_i = \u_issue.slot0_valid_r ? fangyuan360 : _3086_;
  assign \u_csr.opcode_opcode_i = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_fifo.data0_out_o : _3087_;
  assign \u_issue.opcode_b_valid_r = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec1.valid_i : 1'h0;
  assign \u_issue.opcode_a_valid_r = \u_issue.slot0_valid_r ? 1'h1 : _3088_;
  assign _3106_ = _3283_ ? 1'h1 : 1'h0;
  assign _3101_ = _3266_ ? 1'h1 : 1'h0;
  assign _3099_ = _3266_ ? 1'h0 : _3106_;
  assign _3093_ = _3265_ ? 1'h1 : 1'h0;
  assign _3094_ = _3265_ ? 1'h0 : _3101_;
  assign _3083_ = _3265_ ? 1'h0 : _3099_;
  assign \u_issue.slot1_valid_r = _3282_ ? 1'h0 : _3094_;
  assign \u_issue.slot0_valid_r = _3282_ ? 1'h0 : _3093_;
  assign \u_frontend.u_npc.branch_request_i = _3282_ ? 1'h0 : _3083_;
  assign _3412_ = \u_issue.single_issue_w ? _3122_ : \u_issue.pc_x_q ;
  assign _3413_ = \u_issue.dual_issue_w ? _3121_ : _3412_;
  assign _3414_ = \u_exec0.branch_d_request_o ? \u_exec0.branch_target_r : _3413_;
  assign _3415_ = \u_exec1.branch_d_request_o ? \u_exec1.branch_target_r : _3414_;
  assign _3416_ = \u_csr.branch_q ? \u_csr.branch_target_q : _3415_;
  assign _3073_ = rst_i ? 32'h00000000 : _3416_;
  logic [5:0] fangyuan361;
  assign fangyuan361 = { \u_issue.u_pipe0_ctrl.exception_wb_q [0], \u_issue.u_pipe0_ctrl.exception_wb_q [1], \u_issue.u_pipe0_ctrl.exception_wb_q [2], \u_issue.u_pipe0_ctrl.exception_wb_q [3], \u_issue.u_pipe0_ctrl.exception_wb_q [4], \u_issue.u_pipe0_ctrl.exception_wb_q [5] };
  assign _3417_ = | fangyuan361;
  logic [4:0] fangyuan362;
  assign fangyuan362 = { \u_csr.opcode_opcode_i [7], \u_csr.opcode_opcode_i [8], \u_csr.opcode_opcode_i [9], \u_csr.opcode_opcode_i [10], \u_csr.opcode_opcode_i [11] };
  assign _3418_ = | fangyuan362;
  always @(_3112_ or \u_csr.opcode_opcode_i [19:15]) begin
    casez (\u_csr.opcode_opcode_i [19:15])
      0:
        _3419_ = _3112_ [0:0] ;
      1:
        _3419_ = _3112_ [1:1] ;
      2:
        _3419_ = _3112_ [2:2] ;
      3:
        _3419_ = _3112_ [3:3] ;
      4:
        _3419_ = _3112_ [4:4] ;
      5:
        _3419_ = _3112_ [5:5] ;
      6:
        _3419_ = _3112_ [6:6] ;
      7:
        _3419_ = _3112_ [7:7] ;
      8:
        _3419_ = _3112_ [8:8] ;
      9:
        _3419_ = _3112_ [9:9] ;
      10:
        _3419_ = _3112_ [10:10] ;
      11:
        _3419_ = _3112_ [11:11] ;
      12:
        _3419_ = _3112_ [12:12] ;
      13:
        _3419_ = _3112_ [13:13] ;
      14:
        _3419_ = _3112_ [14:14] ;
      15:
        _3419_ = _3112_ [15:15] ;
      16:
        _3419_ = _3112_ [16:16] ;
      17:
        _3419_ = _3112_ [17:17] ;
      18:
        _3419_ = _3112_ [18:18] ;
      19:
        _3419_ = _3112_ [19:19] ;
      20:
        _3419_ = _3112_ [20:20] ;
      21:
        _3419_ = _3112_ [21:21] ;
      22:
        _3419_ = _3112_ [22:22] ;
      23:
        _3419_ = _3112_ [23:23] ;
      24:
        _3419_ = _3112_ [24:24] ;
      25:
        _3419_ = _3112_ [25:25] ;
      26:
        _3419_ = _3112_ [26:26] ;
      27:
        _3419_ = _3112_ [27:27] ;
      28:
        _3419_ = _3112_ [28:28] ;
      29:
        _3419_ = _3112_ [29:29] ;
      30:
        _3419_ = _3112_ [30:30] ;
      31:
        _3419_ = _3112_ [31:31] ;
    endcase
  end
  always @(_3112_ or \u_csr.opcode_opcode_i [24:20]) begin
    casez (\u_csr.opcode_opcode_i [24:20])
      0:
        _3420_ = _3112_ [0:0] ;
      1:
        _3420_ = _3112_ [1:1] ;
      2:
        _3420_ = _3112_ [2:2] ;
      3:
        _3420_ = _3112_ [3:3] ;
      4:
        _3420_ = _3112_ [4:4] ;
      5:
        _3420_ = _3112_ [5:5] ;
      6:
        _3420_ = _3112_ [6:6] ;
      7:
        _3420_ = _3112_ [7:7] ;
      8:
        _3420_ = _3112_ [8:8] ;
      9:
        _3420_ = _3112_ [9:9] ;
      10:
        _3420_ = _3112_ [10:10] ;
      11:
        _3420_ = _3112_ [11:11] ;
      12:
        _3420_ = _3112_ [12:12] ;
      13:
        _3420_ = _3112_ [13:13] ;
      14:
        _3420_ = _3112_ [14:14] ;
      15:
        _3420_ = _3112_ [15:15] ;
      16:
        _3420_ = _3112_ [16:16] ;
      17:
        _3420_ = _3112_ [17:17] ;
      18:
        _3420_ = _3112_ [18:18] ;
      19:
        _3420_ = _3112_ [19:19] ;
      20:
        _3420_ = _3112_ [20:20] ;
      21:
        _3420_ = _3112_ [21:21] ;
      22:
        _3420_ = _3112_ [22:22] ;
      23:
        _3420_ = _3112_ [23:23] ;
      24:
        _3420_ = _3112_ [24:24] ;
      25:
        _3420_ = _3112_ [25:25] ;
      26:
        _3420_ = _3112_ [26:26] ;
      27:
        _3420_ = _3112_ [27:27] ;
      28:
        _3420_ = _3112_ [28:28] ;
      29:
        _3420_ = _3112_ [29:29] ;
      30:
        _3420_ = _3112_ [30:30] ;
      31:
        _3420_ = _3112_ [31:31] ;
    endcase
  end
  always @(_3112_ or \u_csr.opcode_opcode_i [11:7]) begin
    casez (\u_csr.opcode_opcode_i [11:7])
      0:
        _3421_ = _3112_ [0:0] ;
      1:
        _3421_ = _3112_ [1:1] ;
      2:
        _3421_ = _3112_ [2:2] ;
      3:
        _3421_ = _3112_ [3:3] ;
      4:
        _3421_ = _3112_ [4:4] ;
      5:
        _3421_ = _3112_ [5:5] ;
      6:
        _3421_ = _3112_ [6:6] ;
      7:
        _3421_ = _3112_ [7:7] ;
      8:
        _3421_ = _3112_ [8:8] ;
      9:
        _3421_ = _3112_ [9:9] ;
      10:
        _3421_ = _3112_ [10:10] ;
      11:
        _3421_ = _3112_ [11:11] ;
      12:
        _3421_ = _3112_ [12:12] ;
      13:
        _3421_ = _3112_ [13:13] ;
      14:
        _3421_ = _3112_ [14:14] ;
      15:
        _3421_ = _3112_ [15:15] ;
      16:
        _3421_ = _3112_ [16:16] ;
      17:
        _3421_ = _3112_ [17:17] ;
      18:
        _3421_ = _3112_ [18:18] ;
      19:
        _3421_ = _3112_ [19:19] ;
      20:
        _3421_ = _3112_ [20:20] ;
      21:
        _3421_ = _3112_ [21:21] ;
      22:
        _3421_ = _3112_ [22:22] ;
      23:
        _3421_ = _3112_ [23:23] ;
      24:
        _3421_ = _3112_ [24:24] ;
      25:
        _3421_ = _3112_ [25:25] ;
      26:
        _3421_ = _3112_ [26:26] ;
      27:
        _3421_ = _3112_ [27:27] ;
      28:
        _3421_ = _3112_ [28:28] ;
      29:
        _3421_ = _3112_ [29:29] ;
      30:
        _3421_ = _3112_ [30:30] ;
      31:
        _3421_ = _3112_ [31:31] ;
    endcase
  end
  always @(_3117_ or \u_exec1.opcode_opcode_i [19:15]) begin
    casez (\u_exec1.opcode_opcode_i [19:15])
      0:
        _3422_ = _3117_ [0:0] ;
      1:
        _3422_ = _3117_ [1:1] ;
      2:
        _3422_ = _3117_ [2:2] ;
      3:
        _3422_ = _3117_ [3:3] ;
      4:
        _3422_ = _3117_ [4:4] ;
      5:
        _3422_ = _3117_ [5:5] ;
      6:
        _3422_ = _3117_ [6:6] ;
      7:
        _3422_ = _3117_ [7:7] ;
      8:
        _3422_ = _3117_ [8:8] ;
      9:
        _3422_ = _3117_ [9:9] ;
      10:
        _3422_ = _3117_ [10:10] ;
      11:
        _3422_ = _3117_ [11:11] ;
      12:
        _3422_ = _3117_ [12:12] ;
      13:
        _3422_ = _3117_ [13:13] ;
      14:
        _3422_ = _3117_ [14:14] ;
      15:
        _3422_ = _3117_ [15:15] ;
      16:
        _3422_ = _3117_ [16:16] ;
      17:
        _3422_ = _3117_ [17:17] ;
      18:
        _3422_ = _3117_ [18:18] ;
      19:
        _3422_ = _3117_ [19:19] ;
      20:
        _3422_ = _3117_ [20:20] ;
      21:
        _3422_ = _3117_ [21:21] ;
      22:
        _3422_ = _3117_ [22:22] ;
      23:
        _3422_ = _3117_ [23:23] ;
      24:
        _3422_ = _3117_ [24:24] ;
      25:
        _3422_ = _3117_ [25:25] ;
      26:
        _3422_ = _3117_ [26:26] ;
      27:
        _3422_ = _3117_ [27:27] ;
      28:
        _3422_ = _3117_ [28:28] ;
      29:
        _3422_ = _3117_ [29:29] ;
      30:
        _3422_ = _3117_ [30:30] ;
      31:
        _3422_ = _3117_ [31:31] ;
    endcase
  end
  always @(_3117_ or \u_exec1.opcode_opcode_i [24:20]) begin
    casez (\u_exec1.opcode_opcode_i [24:20])
      0:
        _3423_ = _3117_ [0:0] ;
      1:
        _3423_ = _3117_ [1:1] ;
      2:
        _3423_ = _3117_ [2:2] ;
      3:
        _3423_ = _3117_ [3:3] ;
      4:
        _3423_ = _3117_ [4:4] ;
      5:
        _3423_ = _3117_ [5:5] ;
      6:
        _3423_ = _3117_ [6:6] ;
      7:
        _3423_ = _3117_ [7:7] ;
      8:
        _3423_ = _3117_ [8:8] ;
      9:
        _3423_ = _3117_ [9:9] ;
      10:
        _3423_ = _3117_ [10:10] ;
      11:
        _3423_ = _3117_ [11:11] ;
      12:
        _3423_ = _3117_ [12:12] ;
      13:
        _3423_ = _3117_ [13:13] ;
      14:
        _3423_ = _3117_ [14:14] ;
      15:
        _3423_ = _3117_ [15:15] ;
      16:
        _3423_ = _3117_ [16:16] ;
      17:
        _3423_ = _3117_ [17:17] ;
      18:
        _3423_ = _3117_ [18:18] ;
      19:
        _3423_ = _3117_ [19:19] ;
      20:
        _3423_ = _3117_ [20:20] ;
      21:
        _3423_ = _3117_ [21:21] ;
      22:
        _3423_ = _3117_ [22:22] ;
      23:
        _3423_ = _3117_ [23:23] ;
      24:
        _3423_ = _3117_ [24:24] ;
      25:
        _3423_ = _3117_ [25:25] ;
      26:
        _3423_ = _3117_ [26:26] ;
      27:
        _3423_ = _3117_ [27:27] ;
      28:
        _3423_ = _3117_ [28:28] ;
      29:
        _3423_ = _3117_ [29:29] ;
      30:
        _3423_ = _3117_ [30:30] ;
      31:
        _3423_ = _3117_ [31:31] ;
    endcase
  end
  always @(_3117_ or \u_exec1.opcode_opcode_i [11:7]) begin
    casez (\u_exec1.opcode_opcode_i [11:7])
      0:
        _3424_ = _3117_ [0:0] ;
      1:
        _3424_ = _3117_ [1:1] ;
      2:
        _3424_ = _3117_ [2:2] ;
      3:
        _3424_ = _3117_ [3:3] ;
      4:
        _3424_ = _3117_ [4:4] ;
      5:
        _3424_ = _3117_ [5:5] ;
      6:
        _3424_ = _3117_ [6:6] ;
      7:
        _3424_ = _3117_ [7:7] ;
      8:
        _3424_ = _3117_ [8:8] ;
      9:
        _3424_ = _3117_ [9:9] ;
      10:
        _3424_ = _3117_ [10:10] ;
      11:
        _3424_ = _3117_ [11:11] ;
      12:
        _3424_ = _3117_ [12:12] ;
      13:
        _3424_ = _3117_ [13:13] ;
      14:
        _3424_ = _3117_ [14:14] ;
      15:
        _3424_ = _3117_ [15:15] ;
      16:
        _3424_ = _3117_ [16:16] ;
      17:
        _3424_ = _3117_ [17:17] ;
      18:
        _3424_ = _3117_ [18:18] ;
      19:
        _3424_ = _3117_ [19:19] ;
      20:
        _3424_ = _3117_ [20:20] ;
      21:
        _3424_ = _3117_ [21:21] ;
      22:
        _3424_ = _3117_ [22:22] ;
      23:
        _3424_ = _3117_ [23:23] ;
      24:
        _3424_ = _3117_ [24:24] ;
      25:
        _3424_ = _3117_ [25:25] ;
      26:
        _3424_ = _3117_ [26:26] ;
      27:
        _3424_ = _3117_ [27:27] ;
      28:
        _3424_ = _3117_ [28:28] ;
      29:
        _3424_ = _3117_ [29:29] ;
      30:
        _3424_ = _3117_ [30:30] ;
      31:
        _3424_ = _3117_ [31:31] ;
    endcase
  end
  assign \u_frontend.u_fetch.branch_pc_i = \u_csr.branch_q ? \u_csr.branch_target_q : \u_issue.pc_x_q ;
  assign \u_issue.issue_a_sb_alloc_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.rd_valid_o : \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_issue.issue_a_exec_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.exec_o : \u_frontend.u_decode.u_dec1.exec_o ;
  assign \u_issue.issue_a_lsu_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.lsu_o : \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_issue.issue_a_branch_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.branch_o : \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_issue.issue_a_mul_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.mul_o : \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_issue.issue_a_div_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.div_o : \u_frontend.u_decode.u_dec1.div_o ;
  assign \u_issue.issue_a_csr_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.csr_o : \u_frontend.u_decode.u_dec1.csr_o ;
  assign \u_issue.issue_a_invalid_w = \u_issue.slot0_valid_r ? \u_frontend.u_decode.u_dec0.invalid_w : \u_frontend.u_decode.u_dec1.invalid_w ;
  assign _3233_[4:0] = \u_issue.opcode_a_fault_r [1] ? 5'h1c : 5'h00;
  assign \u_issue.issue_a_fault_w = \u_issue.opcode_a_fault_r [0] ? 5'h11 : _3233_[4:0];
  assign _3234_[4:0] = \u_issue.opcode_b_fault_r [1] ? 5'h1c : 5'h00;
  assign \u_issue.issue_b_fault_w = \u_issue.opcode_b_fault_r [0] ? 5'h11 : _3234_[4:0];
  assign \u_csr.u_csrfile.exception_pc_i = _3417_ ? \u_issue.u_pipe0_ctrl.pc_wb_q : \u_issue.u_pipe1_ctrl.pc_wb_q ;
  assign \u_csr.u_csrfile.exception_addr_i = _3417_ ? \u_issue.u_pipe0_ctrl.result_wb_q : \u_issue.u_pipe1_ctrl.result_wb_q ;
  assign \u_frontend.u_npc.branch_source_i = _3133_ ? \u_exec1.pc_m_q : \u_exec0.pc_m_q ;
  assign \u_frontend.u_npc.branch_pc_i = _3133_ ? \u_exec1.pc_x_q : \u_exec0.pc_x_q ;
  assign _3425_ = \u_issue.pipe1_mux_lsu_r ? \u_exec1.opcode_valid_i : \u_div.opcode_valid_i ;
  assign \u_issue.mul_opcode_valid_o = \u_issue.pipe1_mux_mul_r ? \u_exec1.opcode_valid_i : \u_div.opcode_valid_i ;
  assign \u_issue.lsu_opcode_opcode_o = \u_issue.pipe1_mux_lsu_r ? \u_exec1.opcode_opcode_i : \u_csr.opcode_opcode_i ;
  assign \u_issue.lsu_opcode_ra_operand_o = \u_issue.pipe1_mux_lsu_r ? \u_exec1.opcode_ra_operand_i : \u_csr.opcode_ra_operand_i ;
  assign \u_issue.lsu_opcode_rb_operand_o = \u_issue.pipe1_mux_lsu_r ? \u_exec1.opcode_rb_operand_i : \u_div.opcode_rb_operand_i ;
  assign \u_issue.mul_opcode_opcode_o = \u_issue.pipe1_mux_mul_r ? \u_exec1.opcode_opcode_i : \u_csr.opcode_opcode_i ;
  assign \u_issue.mul_opcode_ra_operand_o = \u_issue.pipe1_mux_mul_r ? \u_exec1.opcode_ra_operand_i : \u_csr.opcode_ra_operand_i ;
  assign \u_issue.mul_opcode_rb_operand_o = \u_issue.pipe1_mux_mul_r ? \u_exec1.opcode_rb_operand_i : \u_div.opcode_rb_operand_i ;
  assign _3449_ = \u_issue.issue_a_lsu_w & \u_issue.issue_a_sb_alloc_w ;
  assign _3450_ = _3449_ & _3480_;
  assign _3451_ = \u_issue.issue_a_lsu_w & _3481_;
  assign _3452_ = _3451_ & _3480_;
  assign _3453_ = \u_issue.issue_a_csr_w & _3480_;
  assign _3454_ = \u_issue.issue_a_div_w & _3480_;
  assign _3455_ = \u_issue.issue_a_mul_w & _3480_;
  assign _3456_ = \u_issue.issue_a_branch_w & _3480_;
  assign _3457_ = \u_issue.issue_a_sb_alloc_w & _3480_;
  logic [4:0] fangyuan363;
  assign fangyuan363 = { \u_issue.u_pipe0_ctrl.ctrl_e1_q [7], \u_issue.u_pipe0_ctrl.ctrl_e1_q [7], \u_issue.u_pipe0_ctrl.ctrl_e1_q [7], \u_issue.u_pipe0_ctrl.ctrl_e1_q [7], \u_issue.u_pipe0_ctrl.ctrl_e1_q [7] };
  assign \u_issue.pipe0_rd_e1_w = fangyuan363 & \u_issue.u_pipe0_ctrl.opcode_e1_q [11:7];
  assign \u_issue.u_pipe0_ctrl.valid_e2_w = \u_issue.u_pipe0_ctrl.valid_e2_q & _3482_;
  logic [4:0] fangyuan364;
  assign fangyuan364 = { _3467_, _3467_, _3467_, _3467_, _3467_ };
  assign \u_issue.pipe0_rd_e2_w = fangyuan364 & \u_issue.u_pipe0_ctrl.opcode_e2_q [11:7];
  assign _3458_ = _3489_ & _3485_;
  assign _3459_ = \u_issue.u_pipe0_ctrl.ctrl_e2_q & 10'h37f;
  assign \u_issue.u_pipe0_ctrl.valid_wb_o = \u_issue.u_pipe0_ctrl.valid_wb_q & _3482_;
  assign \u_issue.pipe0_csr_wb_w = \u_issue.u_pipe0_ctrl.ctrl_wb_q [3] & _3482_;
  logic [4:0] fangyuan365;
  assign fangyuan365 = { _3474_, _3474_, _3474_, _3474_, _3474_ };
  assign \u_issue.pipe0_rd_wb_w = fangyuan365 & \u_issue.u_pipe0_ctrl.opcode_wb_q [11:7];
  assign \u_issue.u_pipe0_ctrl.branch_misaligned_w = \u_exec0.branch_d_request_o && _3477_;
  assign _3461_ = \u_div.opcode_valid_i && \u_div.opcode_valid_i ;
  assign _3462_ = _3461_ && _3478_;
  assign _3463_ = $signed(32'h00000001) && \u_issue.u_pipe0_ctrl.valid_e2_w ;
  assign _3464_ = _3463_ && _3476_;
  assign _3465_ = _3463_ && \u_issue.u_pipe0_ctrl.ctrl_e2_q [5];
  assign _3466_ = \u_issue.u_pipe0_ctrl.valid_e2_w && \u_issue.u_pipe0_ctrl.ctrl_e2_q [7];
  assign _3467_ = _3466_ && _3483_;
  assign _3468_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [4] && _3484_;
  assign _3469_ = \u_issue.u_pipe0_ctrl.valid_e2_q && _3476_;
  assign _3470_ = _3469_ && \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign _3471_ = \u_issue.u_pipe0_ctrl.valid_e2_w && _3476_;
  assign _3472_ = \u_issue.u_pipe0_ctrl.valid_e2_w && \u_issue.u_pipe0_ctrl.ctrl_e2_q [5];
  assign _3473_ = \u_issue.u_pipe0_ctrl.valid_wb_o && \u_issue.u_pipe0_ctrl.ctrl_wb_q [7];
  assign _3474_ = _3473_ && _3483_;
  assign _3475_ = \u_issue.pipe0_squash_e1_e2_w || \u_issue.pipe1_squash_e1_e2_w ;
  assign _3476_ = \u_issue.u_pipe0_ctrl.ctrl_e2_q [1] || \u_issue.u_pipe0_ctrl.ctrl_e2_q [2];
  assign \u_issue.pipe0_stall_raw_w = _3468_ || _3458_;
  assign _3477_ = | \u_exec0.branch_target_r [1:0];
  assign _3478_ = ~ _3475_;
  assign _3479_ = ~ _3488_;
  assign _3480_ = ~ \u_csr.take_interrupt_q ;
  assign _3481_ = ~ \u_issue.issue_a_sb_alloc_w ;
  assign _3482_ = ~ \u_exec0.hold_i ;
  assign _3483_ = ~ \u_issue.pipe0_stall_raw_w ;
  assign _3484_ = ~ \u_div.valid_q ;
  assign _3485_ = ~ \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign _3486_ = \u_issue.issue_a_lsu_w | \u_issue.issue_a_csr_w ;
  assign _3487_ = _3486_ | \u_issue.issue_a_div_w ;
  assign _3488_ = _3487_ | \u_issue.issue_a_mul_w ;
  assign _3489_ = \u_issue.u_pipe0_ctrl.ctrl_e2_q [1] | \u_issue.u_pipe0_ctrl.ctrl_e2_q [2];
  assign \u_issue.pipe0_squash_e1_e2_w = \u_issue.u_pipe0_ctrl.squash_e1_e2_w | \u_issue.u_pipe0_ctrl.squash_e1_e2_q ;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.valid_wb_q <= _3447_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.ctrl_wb_q <= _3432_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.csr_wr_wb_q <= _3429_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.csr_wdata_wb_q <= _3427_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.result_wb_q <= _3443_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.pc_wb_q <= _3441_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.opcode_wb_q <= _3438_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.exception_wb_q <= _3435_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.squash_e1_e2_q <= _3444_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.result_e2_q <= _3442_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.valid_e2_q <= _3446_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.ctrl_e2_q <= _3431_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.csr_wr_e2_q <= _3428_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.csr_wdata_e2_q <= _3426_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.pc_e2_q <= _3440_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.opcode_e2_q <= _3437_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.exception_e2_q <= _3434_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.exception_e1_q <= _3433_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.valid_e1_q <= _3445_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.ctrl_e1_q <= _3430_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.pc_e1_q <= _3439_;
  always @(posedge clk_i)
      \u_issue.u_pipe0_ctrl.opcode_e1_q <= _3436_;
  assign _3490_ = 1'h0 ? 6'h00 : \u_issue.u_pipe0_ctrl.exception_e2_r ;
  assign _3491_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.exception_wb_q : _3490_;
  assign _3435_ = rst_i ? 6'h00 : _3491_;
  assign _3492_ = 1'h0 ? 32'h00000000 : \u_issue.u_pipe0_ctrl.opcode_e2_q ;
  assign _3493_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.opcode_wb_q : _3492_;
  assign _3438_ = rst_i ? 32'h00000000 : _3493_;
  assign _3494_ = 1'h0 ? 32'h00000000 : \u_issue.u_pipe0_ctrl.pc_e2_q ;
  assign _3495_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.pc_wb_q : _3494_;
  assign _3441_ = rst_i ? 32'h00000000 : _3495_;
  assign _3496_ = _3472_ ? \u_mul.result_e2_q : \u_issue.u_pipe0_ctrl.result_e2_q ;
  assign _3497_ = _3471_ ? \u_issue.u_pipe0_ctrl.mem_result_e2_i : _3496_;
  assign _3498_ = 1'h0 ? 32'h00000000 : _3497_;
  assign _3499_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.result_wb_q : _3498_;
  assign _3443_ = rst_i ? 32'h00000000 : _3499_;
  assign _3500_ = 1'h0 ? 32'h00000000 : \u_issue.u_pipe0_ctrl.csr_wdata_e2_q ;
  assign _3501_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.csr_wdata_wb_q : _3500_;
  assign _3427_ = rst_i ? 32'h00000000 : _3501_;
  assign _3502_ = 1'h0 ? 1'h0 : \u_issue.u_pipe0_ctrl.csr_wr_e2_q ;
  assign _3503_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.csr_wr_wb_q : _3502_;
  assign _3429_ = rst_i ? 1'h0 : _3503_;
  assign _3504_ = \u_issue.u_pipe0_ctrl.squash_e1_e2_w ? _3459_ : \u_issue.u_pipe0_ctrl.ctrl_e2_q ;
  assign _3505_ = 1'h0 ? 10'h000 : _3504_;
  assign _3506_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_wb_q : _3505_;
  assign _3432_ = rst_i ? 10'h000 : _3506_;
  assign _3507_ = _3509_ ? 1'h0 : \u_issue.u_pipe0_ctrl.valid_e2_q ;
  logic [5:0] fangyuan366;
  assign fangyuan366 = { _3508_[0], _3508_[1], _3508_[2], _3508_[3], _3508_[4], _3508_[5] };
  assign _3509_ = | fangyuan366;
  assign _3508_[0] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h14;
  assign _3508_[1] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h15;
  assign _3508_[2] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h16;
  assign _3508_[3] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h17;
  assign _3508_[4] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h1d;
  assign _3508_[5] = \u_issue.u_pipe0_ctrl.exception_e2_r == 5'h1f;
  assign _3510_ = 1'h0 ? 1'h0 : _3507_;
  assign _3511_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.valid_wb_q : _3510_;
  assign _3447_ = rst_i ? 1'h0 : _3511_;
  assign _3512_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.squash_e1_e2_q : \u_issue.u_pipe0_ctrl.squash_e1_e2_w ;
  assign _3444_ = rst_i ? 1'h0 : _3512_;
  logic [5:0] fangyuan367;
  assign fangyuan367 = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign \u_issue.u_pipe0_ctrl.exception_e2_r = _3470_ ? fangyuan367 : \u_issue.u_pipe0_ctrl.exception_e2_q ;
  assign _3448_ = _3465_ ? \u_mul.result_e2_q : \u_issue.u_pipe0_ctrl.result_e2_q ;
  assign \u_issue.pipe0_result_e2_w = _3464_ ? \u_issue.u_pipe0_ctrl.mem_result_e2_i : _3448_;
  assign _3513_ = _3514_ ? \u_issue.u_pipe0_ctrl.exception_e1_q : \u_csr.exception_e1_q ;
  assign _3515_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [8] ? 6'h20 : _3513_;
  assign _3516_ = _3475_ ? 6'h00 : _3515_;
  assign _3517_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.exception_e2_q : _3516_;
  assign _3434_ = rst_i ? 6'h00 : _3517_;
  assign _3518_ = _3475_ ? 32'h00000000 : \u_issue.u_pipe0_ctrl.opcode_e1_q ;
  assign _3519_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.opcode_e2_q : _3518_;
  assign _3437_ = rst_i ? 32'h00000000 : _3519_;
  assign _3520_ = _3475_ ? 32'h00000000 : \u_issue.u_pipe0_ctrl.pc_e1_q ;
  assign _3521_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.pc_e2_q : _3520_;
  assign _3440_ = rst_i ? 32'h00000000 : _3521_;
  assign _3522_ = _3475_ ? 32'h00000000 : \u_csr.csr_wdata_e1_q ;
  assign _3523_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.csr_wdata_e2_q : _3522_;
  assign _3426_ = rst_i ? 32'h00000000 : _3523_;
  assign _3524_ = _3475_ ? 1'h0 : \u_csr.rd_valid_e1_q ;
  assign _3525_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.csr_wr_e2_q : _3524_;
  assign _3428_ = rst_i ? 1'h0 : _3525_;
  assign _3526_ = _3475_ ? 10'h000 : \u_issue.u_pipe0_ctrl.ctrl_e1_q ;
  assign _3527_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e2_q : _3526_;
  assign _3431_ = rst_i ? 10'h000 : _3527_;
  assign _3528_ = _3514_ ? 1'h0 : \u_issue.u_pipe0_ctrl.valid_e1_q ;
  assign _3529_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [8] ? \u_issue.u_pipe0_ctrl.valid_e1_q : _3528_;
  assign _3530_ = _3475_ ? 1'h0 : _3529_;
  assign _3531_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.valid_e2_q : _3530_;
  assign _3446_ = rst_i ? 1'h0 : _3531_;
  assign _3532_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [3] ? \u_csr.rd_result_e1_q : \u_exec0.result_q ;
  assign _3533_ = \u_issue.u_pipe0_ctrl.ctrl_e1_q [4] ? \u_div.wb_result_q : _3532_;
  assign _3534_ = _3475_ ? 32'h00000000 : _3533_;
  assign _3535_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.result_e2_q : _3534_;
  assign _3442_ = rst_i ? 32'h00000000 : _3535_;
  assign _3536_ = _3462_ ? 1'h1 : 1'h0;
  assign _3537_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [9] : _3536_;
  assign _3430_[9] = rst_i ? 1'h0 : _3537_;
  assign _3538_ = _3462_ ? _3457_ : 1'h0;
  assign _3539_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [7] : _3538_;
  assign _3430_[7] = rst_i ? 1'h0 : _3539_;
  assign _3540_ = _3462_ ? _3456_ : 1'h0;
  assign _3541_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [6] : _3540_;
  assign _3430_[6] = rst_i ? 1'h0 : _3541_;
  assign _3542_ = _3462_ ? _3455_ : 1'h0;
  assign _3543_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [5] : _3542_;
  assign _3430_[5] = rst_i ? 1'h0 : _3543_;
  assign _3544_ = _3462_ ? _3454_ : 1'h0;
  assign _3545_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [4] : _3544_;
  assign _3430_[4] = rst_i ? 1'h0 : _3545_;
  assign _3546_ = _3462_ ? _3453_ : 1'h0;
  assign _3547_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [3] : _3546_;
  assign _3430_[3] = rst_i ? 1'h0 : _3547_;
  assign _3548_ = _3462_ ? _3452_ : 1'h0;
  assign _3549_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [2] : _3548_;
  assign _3430_[2] = rst_i ? 1'h0 : _3549_;
  assign _3550_ = _3462_ ? _3450_ : 1'h0;
  assign _3551_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [1] : _3550_;
  assign _3430_[1] = rst_i ? 1'h0 : _3551_;
  assign _3552_ = _3462_ ? _3479_ : 1'h0;
  assign _3553_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [0] : _3552_;
  assign _3430_[0] = rst_i ? 1'h0 : _3553_;
  assign _3554_ = _3462_ ? \u_csr.take_interrupt_q : 1'h0;
  assign _3555_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.ctrl_e1_q [8] : _3554_;
  assign _3430_[8] = rst_i ? 1'h0 : _3555_;
  assign _3556_ = _3462_ ? \u_csr.opcode_opcode_i : 32'h00000000;
  assign _3557_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.opcode_e1_q : _3556_;
  assign _3436_ = rst_i ? 32'h00000000 : _3557_;
  assign _3558_ = _3462_ ? \u_exec0.opcode_pc_i : 32'h00000000;
  assign _3559_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.pc_e1_q : _3558_;
  assign _3439_ = rst_i ? 32'h00000000 : _3559_;
  assign _3560_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.valid_e1_q : _3536_;
  assign _3445_ = rst_i ? 1'h0 : _3560_;
  assign _3561_ = _3462_ ? _3564_ : 6'h00;
  assign _3562_ = \u_exec0.hold_i ? \u_issue.u_pipe0_ctrl.exception_e1_q : _3561_;
  assign _3433_ = rst_i ? 6'h00 : _3562_;
  logic [5:0] fangyuan368;
  assign fangyuan368 = { \u_issue.issue_a_fault_w [0], \u_issue.issue_a_fault_w [1], \u_issue.issue_a_fault_w [2], \u_issue.issue_a_fault_w [3], \u_issue.issue_a_fault_w [4], 1'h0 };
  assign _3563_ = | fangyuan368;
  logic [5:0] fangyuan369;
  assign fangyuan369 = { \u_issue.u_pipe0_ctrl.exception_e1_q [0], \u_issue.u_pipe0_ctrl.exception_e1_q [1], \u_issue.u_pipe0_ctrl.exception_e1_q [2], \u_issue.u_pipe0_ctrl.exception_e1_q [3], \u_issue.u_pipe0_ctrl.exception_e1_q [4], \u_issue.u_pipe0_ctrl.exception_e1_q [5] };
  assign _3514_ = | fangyuan369;
  logic [5:0] fangyuan370;
  assign fangyuan370 = { \u_issue.u_pipe0_ctrl.exception_e2_r [0], \u_issue.u_pipe0_ctrl.exception_e2_r [1], \u_issue.u_pipe0_ctrl.exception_e2_r [2], \u_issue.u_pipe0_ctrl.exception_e2_r [3], \u_issue.u_pipe0_ctrl.exception_e2_r [4], \u_issue.u_pipe0_ctrl.exception_e2_r [5] };
  assign \u_issue.u_pipe0_ctrl.squash_e1_e2_w = | fangyuan370;
  assign _3460_[4:0] = \u_issue.u_pipe0_ctrl.branch_misaligned_w ? 5'h10 : 5'h00;
  logic [5:0] fangyuan371;
  assign fangyuan371 = { 1'h0, \u_issue.issue_a_fault_w };
  logic [5:0] fangyuan372;
  assign fangyuan372 = { 1'h0, _3460_[4:0] };
  assign _3564_ = _3563_ ? fangyuan371 : fangyuan372;
  assign _3584_ = \u_frontend.u_decode.u_dec1.lsu_o & \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign _3585_ = _3584_ & _3615_;
  assign _3586_ = \u_frontend.u_decode.u_dec1.lsu_o & _3616_;
  assign _3587_ = _3586_ & _3615_;
  assign _3588_ = 1'h0 & _3615_;
  assign _3589_ = 1'h0 & _3615_;
  assign _3590_ = \u_frontend.u_decode.u_dec1.mul_o & _3615_;
  assign _3591_ = \u_frontend.u_decode.u_dec1.branch_o & _3615_;
  assign _3592_ = \u_frontend.u_decode.u_dec1.rd_valid_o & _3615_;
  logic [4:0] fangyuan373;
  assign fangyuan373 = { \u_issue.u_pipe1_ctrl.ctrl_e1_q [7], \u_issue.u_pipe1_ctrl.ctrl_e1_q [7], \u_issue.u_pipe1_ctrl.ctrl_e1_q [7], \u_issue.u_pipe1_ctrl.ctrl_e1_q [7], \u_issue.u_pipe1_ctrl.ctrl_e1_q [7] };
  assign \u_issue.pipe1_rd_e1_w = fangyuan373 & \u_issue.u_pipe1_ctrl.opcode_e1_q [11:7];
  assign \u_issue.u_pipe1_ctrl.valid_e2_w = \u_issue.u_pipe1_ctrl.valid_e2_q & _3617_;
  logic [4:0] fangyuan374;
  assign fangyuan374 = { _3602_, _3602_, _3602_, _3602_, _3602_ };
  assign \u_issue.pipe1_rd_e2_w = fangyuan374 & \u_issue.u_pipe1_ctrl.opcode_e2_q [11:7];
  assign _3593_ = _3624_ & _3620_;
  assign _3594_ = \u_issue.u_pipe1_ctrl.ctrl_e2_q & 10'h37f;
  assign \u_issue.u_pipe1_ctrl.valid_wb_o = \u_issue.u_pipe1_ctrl.valid_wb_q & _3617_;
  logic [4:0] fangyuan375;
  assign fangyuan375 = { _3609_, _3609_, _3609_, _3609_, _3609_ };
  assign \u_issue.pipe1_rd_wb_w = fangyuan375 & \u_issue.u_pipe1_ctrl.opcode_wb_q [11:7];
  assign \u_issue.u_pipe1_ctrl.branch_misaligned_w = \u_exec1.branch_d_request_o && _3612_;
  assign _3596_ = \u_exec1.opcode_valid_i && \u_exec1.opcode_valid_i ;
  assign _3597_ = _3596_ && _3613_;
  assign _3598_ = $signed(32'h00000001) && \u_issue.u_pipe1_ctrl.valid_e2_w ;
  assign _3599_ = _3598_ && _3611_;
  assign _3600_ = _3598_ && \u_issue.u_pipe1_ctrl.ctrl_e2_q [5];
  assign _3601_ = \u_issue.u_pipe1_ctrl.valid_e2_w && \u_issue.u_pipe1_ctrl.ctrl_e2_q [7];
  assign _3602_ = _3601_ && _3618_;
  assign _3603_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [4] && _3619_;
  assign _3604_ = \u_issue.u_pipe1_ctrl.valid_e2_q && _3611_;
  assign _3605_ = _3604_ && \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign _3606_ = \u_issue.u_pipe1_ctrl.valid_e2_w && _3611_;
  assign _3607_ = \u_issue.u_pipe1_ctrl.valid_e2_w && \u_issue.u_pipe1_ctrl.ctrl_e2_q [5];
  assign _3608_ = \u_issue.u_pipe1_ctrl.valid_wb_o && \u_issue.u_pipe1_ctrl.ctrl_wb_q [7];
  assign _3609_ = _3608_ && _3618_;
  assign _3610_ = \u_issue.pipe1_squash_e1_e2_w || \u_issue.pipe0_squash_e1_e2_w ;
  assign _3611_ = \u_issue.u_pipe1_ctrl.ctrl_e2_q [1] || \u_issue.u_pipe1_ctrl.ctrl_e2_q [2];
  assign \u_issue.pipe1_stall_raw_w = _3603_ || _3593_;
  assign _3612_ = | \u_exec1.branch_target_r [1:0];
  assign _3613_ = ~ _3610_;
  assign _3614_ = ~ _3623_;
  assign _3615_ = ~ \u_csr.take_interrupt_q ;
  assign _3616_ = ~ \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign _3617_ = ~ \u_exec0.hold_i ;
  assign _3618_ = ~ \u_issue.pipe1_stall_raw_w ;
  assign _3619_ = ~ \u_div.valid_q ;
  assign _3620_ = ~ \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign _3621_ = \u_frontend.u_decode.u_dec1.lsu_o | 1'h0;
  assign _3622_ = _3621_ | 1'h0;
  assign _3623_ = _3622_ | \u_frontend.u_decode.u_dec1.mul_o ;
  assign _3624_ = \u_issue.u_pipe1_ctrl.ctrl_e2_q [1] | \u_issue.u_pipe1_ctrl.ctrl_e2_q [2];
  assign \u_issue.pipe1_squash_e1_e2_w = \u_issue.u_pipe1_ctrl.squash_e1_e2_w | \u_issue.u_pipe1_ctrl.squash_e1_e2_q ;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.valid_wb_q <= _3582_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.ctrl_wb_q <= _3567_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.result_wb_q <= _3578_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.pc_wb_q <= _3576_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.opcode_wb_q <= _3573_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.exception_wb_q <= _3570_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.squash_e1_e2_q <= _3579_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.result_e2_q <= _3577_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.valid_e2_q <= _3581_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.ctrl_e2_q <= _3566_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.pc_e2_q <= _3575_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.opcode_e2_q <= _3572_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.exception_e2_q <= _3569_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.exception_e1_q <= _3568_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.valid_e1_q <= _3580_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.ctrl_e1_q <= _3565_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.pc_e1_q <= _3574_;
  always @(posedge clk_i)
      \u_issue.u_pipe1_ctrl.opcode_e1_q <= _3571_;
  assign _3625_ = \u_issue.pipe0_squash_e1_e2_w ? 6'h00 : \u_issue.u_pipe1_ctrl.exception_e2_r ;
  assign _3626_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.exception_wb_q : _3625_;
  assign _3570_ = rst_i ? 6'h00 : _3626_;
  assign _3627_ = \u_issue.pipe0_squash_e1_e2_w ? 32'h00000000 : \u_issue.u_pipe1_ctrl.opcode_e2_q ;
  assign _3628_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.opcode_wb_q : _3627_;
  assign _3573_ = rst_i ? 32'h00000000 : _3628_;
  assign _3629_ = \u_issue.pipe0_squash_e1_e2_w ? 32'h00000000 : \u_issue.u_pipe1_ctrl.pc_e2_q ;
  assign _3630_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.pc_wb_q : _3629_;
  assign _3576_ = rst_i ? 32'h00000000 : _3630_;
  assign _3631_ = _3607_ ? \u_mul.result_e2_q : \u_issue.u_pipe1_ctrl.result_e2_q ;
  assign _3632_ = _3606_ ? \u_issue.u_pipe0_ctrl.mem_result_e2_i : _3631_;
  assign _3633_ = \u_issue.pipe0_squash_e1_e2_w ? 32'h00000000 : _3632_;
  assign _3634_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.result_wb_q : _3633_;
  assign _3578_ = rst_i ? 32'h00000000 : _3634_;
  assign _3635_ = \u_issue.u_pipe1_ctrl.squash_e1_e2_w ? _3594_ : \u_issue.u_pipe1_ctrl.ctrl_e2_q ;
  assign _3636_ = \u_issue.pipe0_squash_e1_e2_w ? 10'h000 : _3635_;
  assign _3637_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_wb_q : _3636_;
  assign _3567_ = rst_i ? 10'h000 : _3637_;
  assign _3638_ = _3640_ ? 1'h0 : \u_issue.u_pipe1_ctrl.valid_e2_q ;
  logic [5:0] fangyuan376;
  assign fangyuan376 = { _3639_[0], _3639_[1], _3639_[2], _3639_[3], _3639_[4], _3639_[5] };
  assign _3640_ = | fangyuan376;
  assign _3639_[0] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h14;
  assign _3639_[1] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h15;
  assign _3639_[2] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h16;
  assign _3639_[3] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h17;
  assign _3639_[4] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h1d;
  assign _3639_[5] = \u_issue.u_pipe1_ctrl.exception_e2_r == 5'h1f;
  assign _3641_ = \u_issue.pipe0_squash_e1_e2_w ? 1'h0 : _3638_;
  assign _3642_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.valid_wb_q : _3641_;
  assign _3582_ = rst_i ? 1'h0 : _3642_;
  assign _3643_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.squash_e1_e2_q : \u_issue.u_pipe1_ctrl.squash_e1_e2_w ;
  assign _3579_ = rst_i ? 1'h0 : _3643_;
  logic [5:0] fangyuan377;
  assign fangyuan377 = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign \u_issue.u_pipe1_ctrl.exception_e2_r = _3605_ ? fangyuan377 : \u_issue.u_pipe1_ctrl.exception_e2_q ;
  assign _3583_ = _3600_ ? \u_mul.result_e2_q : \u_issue.u_pipe1_ctrl.result_e2_q ;
  assign \u_issue.pipe1_result_e2_w = _3599_ ? \u_issue.u_pipe0_ctrl.mem_result_e2_i : _3583_;
  assign _3644_ = _3645_ ? \u_issue.u_pipe1_ctrl.exception_e1_q : \u_csr.exception_e1_q ;
  assign _3646_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [8] ? 6'h20 : _3644_;
  assign _3647_ = _3610_ ? 6'h00 : _3646_;
  assign _3648_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.exception_e2_q : _3647_;
  assign _3569_ = rst_i ? 6'h00 : _3648_;
  assign _3649_ = _3610_ ? 32'h00000000 : \u_issue.u_pipe1_ctrl.opcode_e1_q ;
  assign _3650_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.opcode_e2_q : _3649_;
  assign _3572_ = rst_i ? 32'h00000000 : _3650_;
  assign _3651_ = _3610_ ? 32'h00000000 : \u_issue.u_pipe1_ctrl.pc_e1_q ;
  assign _3652_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.pc_e2_q : _3651_;
  assign _3575_ = rst_i ? 32'h00000000 : _3652_;
  assign _3653_ = _3610_ ? 10'h000 : \u_issue.u_pipe1_ctrl.ctrl_e1_q ;
  assign _3654_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e2_q : _3653_;
  assign _3566_ = rst_i ? 10'h000 : _3654_;
  assign _3655_ = _3645_ ? 1'h0 : \u_issue.u_pipe1_ctrl.valid_e1_q ;
  assign _3656_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [8] ? \u_issue.u_pipe1_ctrl.valid_e1_q : _3655_;
  assign _3657_ = _3610_ ? 1'h0 : _3656_;
  assign _3658_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.valid_e2_q : _3657_;
  assign _3581_ = rst_i ? 1'h0 : _3658_;
  assign _3659_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [3] ? \u_csr.rd_result_e1_q : \u_exec1.result_q ;
  assign _3660_ = \u_issue.u_pipe1_ctrl.ctrl_e1_q [4] ? \u_div.wb_result_q : _3659_;
  assign _3661_ = _3610_ ? 32'h00000000 : _3660_;
  assign _3662_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.result_e2_q : _3661_;
  assign _3577_ = rst_i ? 32'h00000000 : _3662_;
  assign _3663_ = _3597_ ? 1'h1 : 1'h0;
  assign _3664_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [9] : _3663_;
  assign _3565_[9] = rst_i ? 1'h0 : _3664_;
  assign _3665_ = _3597_ ? _3592_ : 1'h0;
  assign _3666_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [7] : _3665_;
  assign _3565_[7] = rst_i ? 1'h0 : _3666_;
  assign _3667_ = _3597_ ? _3591_ : 1'h0;
  assign _3668_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [6] : _3667_;
  assign _3565_[6] = rst_i ? 1'h0 : _3668_;
  assign _3669_ = _3597_ ? _3590_ : 1'h0;
  assign _3670_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [5] : _3669_;
  assign _3565_[5] = rst_i ? 1'h0 : _3670_;
  assign _3671_ = _3597_ ? _3589_ : 1'h0;
  assign _3672_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [4] : _3671_;
  assign _3565_[4] = rst_i ? 1'h0 : _3672_;
  assign _3673_ = _3597_ ? _3588_ : 1'h0;
  assign _3674_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [3] : _3673_;
  assign _3565_[3] = rst_i ? 1'h0 : _3674_;
  assign _3675_ = _3597_ ? _3587_ : 1'h0;
  assign _3676_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [2] : _3675_;
  assign _3565_[2] = rst_i ? 1'h0 : _3676_;
  assign _3677_ = _3597_ ? _3585_ : 1'h0;
  assign _3678_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [1] : _3677_;
  assign _3565_[1] = rst_i ? 1'h0 : _3678_;
  assign _3679_ = _3597_ ? _3614_ : 1'h0;
  assign _3680_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [0] : _3679_;
  assign _3565_[0] = rst_i ? 1'h0 : _3680_;
  assign _3681_ = _3597_ ? \u_csr.take_interrupt_q : 1'h0;
  assign _3682_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.ctrl_e1_q [8] : _3681_;
  assign _3565_[8] = rst_i ? 1'h0 : _3682_;
  assign _3683_ = _3597_ ? \u_exec1.opcode_opcode_i : 32'h00000000;
  assign _3684_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.opcode_e1_q : _3683_;
  assign _3571_ = rst_i ? 32'h00000000 : _3684_;
  assign _3685_ = _3597_ ? \u_exec1.opcode_pc_i : 32'h00000000;
  assign _3686_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.pc_e1_q : _3685_;
  assign _3574_ = rst_i ? 32'h00000000 : _3686_;
  assign _3687_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.valid_e1_q : _3663_;
  assign _3580_ = rst_i ? 1'h0 : _3687_;
  assign _3688_ = _3597_ ? _3691_ : 6'h00;
  assign _3689_ = \u_exec0.hold_i ? \u_issue.u_pipe1_ctrl.exception_e1_q : _3688_;
  assign _3568_ = rst_i ? 6'h00 : _3689_;
  logic [5:0] fangyuan378;
  assign fangyuan378 = { \u_issue.issue_b_fault_w [0], \u_issue.issue_b_fault_w [1], \u_issue.issue_b_fault_w [2], \u_issue.issue_b_fault_w [3], \u_issue.issue_b_fault_w [4], 1'h0 };
  assign _3690_ = | fangyuan378;
  logic [5:0] fangyuan379;
  assign fangyuan379 = { \u_issue.u_pipe1_ctrl.exception_e1_q [0], \u_issue.u_pipe1_ctrl.exception_e1_q [1], \u_issue.u_pipe1_ctrl.exception_e1_q [2], \u_issue.u_pipe1_ctrl.exception_e1_q [3], \u_issue.u_pipe1_ctrl.exception_e1_q [4], \u_issue.u_pipe1_ctrl.exception_e1_q [5] };
  assign _3645_ = | fangyuan379;
  logic [5:0] fangyuan380;
  assign fangyuan380 = { \u_issue.u_pipe1_ctrl.exception_e2_r [0], \u_issue.u_pipe1_ctrl.exception_e2_r [1], \u_issue.u_pipe1_ctrl.exception_e2_r [2], \u_issue.u_pipe1_ctrl.exception_e2_r [3], \u_issue.u_pipe1_ctrl.exception_e2_r [4], \u_issue.u_pipe1_ctrl.exception_e2_r [5] };
  assign \u_issue.u_pipe1_ctrl.squash_e1_e2_w = | fangyuan380;
  assign _3595_[4:0] = \u_issue.u_pipe1_ctrl.branch_misaligned_w ? 5'h10 : 5'h00;
  logic [5:0] fangyuan381;
  assign fangyuan381 = { 1'h0, \u_issue.issue_b_fault_w };
  logic [5:0] fangyuan382;
  assign fangyuan382 = { 1'h0, _3595_[4:0] };
  assign _3691_ = _3690_ ? fangyuan381 : fangyuan382;
  assign _3723_ = \u_issue.pipe0_rd_wb_w == 1'h1;
  assign _3724_ = \u_issue.pipe1_rd_wb_w == 1'h1;
  assign _3725_ = \u_issue.pipe0_rd_wb_w == 2'h2;
  assign _3726_ = \u_issue.pipe1_rd_wb_w == 2'h2;
  assign _3727_ = \u_issue.pipe0_rd_wb_w == 2'h3;
  assign _3728_ = \u_issue.pipe1_rd_wb_w == 2'h3;
  assign _3729_ = \u_issue.pipe0_rd_wb_w == 3'h4;
  assign _3730_ = \u_issue.pipe1_rd_wb_w == 3'h4;
  assign _3731_ = \u_issue.pipe0_rd_wb_w == 3'h5;
  assign _3732_ = \u_issue.pipe1_rd_wb_w == 3'h5;
  assign _3733_ = \u_issue.pipe0_rd_wb_w == 3'h6;
  assign _3734_ = \u_issue.pipe1_rd_wb_w == 3'h6;
  assign _3735_ = \u_issue.pipe0_rd_wb_w == 3'h7;
  assign _3736_ = \u_issue.pipe1_rd_wb_w == 3'h7;
  assign _3737_ = \u_issue.pipe0_rd_wb_w == 4'h8;
  assign _3738_ = \u_issue.pipe1_rd_wb_w == 4'h8;
  assign _3739_ = \u_issue.pipe0_rd_wb_w == 4'h9;
  assign _3740_ = \u_issue.pipe1_rd_wb_w == 4'h9;
  assign _3741_ = \u_issue.pipe0_rd_wb_w == 4'ha;
  assign _3742_ = \u_issue.pipe1_rd_wb_w == 4'ha;
  assign _3743_ = \u_issue.pipe0_rd_wb_w == 4'hb;
  assign _3744_ = \u_issue.pipe1_rd_wb_w == 4'hb;
  assign _3745_ = \u_issue.pipe0_rd_wb_w == 4'hc;
  assign _3746_ = \u_issue.pipe1_rd_wb_w == 4'hc;
  assign _3747_ = \u_issue.pipe0_rd_wb_w == 4'hd;
  assign _3748_ = \u_issue.pipe1_rd_wb_w == 4'hd;
  assign _3749_ = \u_issue.pipe0_rd_wb_w == 4'he;
  assign _3750_ = \u_issue.pipe1_rd_wb_w == 4'he;
  assign _3751_ = \u_issue.pipe0_rd_wb_w == 4'hf;
  assign _3752_ = \u_issue.pipe1_rd_wb_w == 4'hf;
  assign _3753_ = \u_issue.pipe0_rd_wb_w == 5'h10;
  assign _3754_ = \u_issue.pipe1_rd_wb_w == 5'h10;
  assign _3755_ = \u_issue.pipe0_rd_wb_w == 5'h11;
  assign _3756_ = \u_issue.pipe1_rd_wb_w == 5'h11;
  assign _3757_ = \u_issue.pipe0_rd_wb_w == 5'h12;
  assign _3758_ = \u_issue.pipe1_rd_wb_w == 5'h12;
  assign _3759_ = \u_issue.pipe0_rd_wb_w == 5'h13;
  assign _3760_ = \u_issue.pipe1_rd_wb_w == 5'h13;
  assign _3761_ = \u_issue.pipe0_rd_wb_w == 5'h14;
  assign _3762_ = \u_issue.pipe1_rd_wb_w == 5'h14;
  assign _3763_ = \u_issue.pipe0_rd_wb_w == 5'h15;
  assign _3764_ = \u_issue.pipe1_rd_wb_w == 5'h15;
  assign _3765_ = \u_issue.pipe0_rd_wb_w == 5'h16;
  assign _3766_ = \u_issue.pipe1_rd_wb_w == 5'h16;
  assign _3767_ = \u_issue.pipe0_rd_wb_w == 5'h17;
  assign _3768_ = \u_issue.pipe1_rd_wb_w == 5'h17;
  assign _3769_ = \u_issue.pipe0_rd_wb_w == 5'h18;
  assign _3770_ = \u_issue.pipe1_rd_wb_w == 5'h18;
  assign _3771_ = \u_issue.pipe0_rd_wb_w == 5'h19;
  assign _3772_ = \u_issue.pipe1_rd_wb_w == 5'h19;
  assign _3773_ = \u_issue.pipe0_rd_wb_w == 5'h1a;
  assign _3774_ = \u_issue.pipe1_rd_wb_w == 5'h1a;
  assign _3775_ = \u_issue.pipe0_rd_wb_w == 5'h1b;
  assign _3776_ = \u_issue.pipe1_rd_wb_w == 5'h1b;
  assign _3777_ = \u_issue.pipe0_rd_wb_w == 5'h1c;
  assign _3778_ = \u_issue.pipe1_rd_wb_w == 5'h1c;
  assign _3779_ = \u_issue.pipe0_rd_wb_w == 5'h1d;
  assign _3780_ = \u_issue.pipe1_rd_wb_w == 5'h1d;
  assign _3781_ = \u_issue.pipe0_rd_wb_w == 5'h1e;
  assign _3782_ = \u_issue.pipe1_rd_wb_w == 5'h1e;
  assign _3783_ = \u_issue.pipe0_rd_wb_w == 5'h1f;
  assign _3784_ = \u_issue.pipe1_rd_wb_w == 5'h1f;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r1_q <= _3702_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r2_q <= _3713_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r3_q <= _3716_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r4_q <= _3717_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r5_q <= _3718_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r6_q <= _3719_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r7_q <= _3720_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r8_q <= _3721_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r9_q <= _3722_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r10_q <= _3692_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r11_q <= _3693_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r12_q <= _3694_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r13_q <= _3695_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r14_q <= _3696_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r15_q <= _3697_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r16_q <= _3698_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r17_q <= _3699_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r18_q <= _3700_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r19_q <= _3701_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r20_q <= _3703_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r21_q <= _3704_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r22_q <= _3705_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r23_q <= _3706_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r24_q <= _3707_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r25_q <= _3708_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r26_q <= _3709_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r27_q <= _3710_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r28_q <= _3711_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r29_q <= _3712_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r30_q <= _3714_;
  always @(posedge clk_i)
      \u_issue.u_regfile.REGFILE.reg_r31_q <= _3715_;
  logic [991:0] fangyuan383;
  assign fangyuan383 = { \u_issue.u_regfile.REGFILE.reg_r1_q , \u_issue.u_regfile.REGFILE.reg_r2_q , \u_issue.u_regfile.REGFILE.reg_r3_q , \u_issue.u_regfile.REGFILE.reg_r4_q , \u_issue.u_regfile.REGFILE.reg_r5_q , \u_issue.u_regfile.REGFILE.reg_r6_q , \u_issue.u_regfile.REGFILE.reg_r7_q , \u_issue.u_regfile.REGFILE.reg_r8_q , \u_issue.u_regfile.REGFILE.reg_r9_q , \u_issue.u_regfile.REGFILE.reg_r10_q , \u_issue.u_regfile.REGFILE.reg_r11_q , \u_issue.u_regfile.REGFILE.reg_r12_q , \u_issue.u_regfile.REGFILE.reg_r13_q , \u_issue.u_regfile.REGFILE.reg_r14_q , \u_issue.u_regfile.REGFILE.reg_r15_q , \u_issue.u_regfile.REGFILE.reg_r16_q , \u_issue.u_regfile.REGFILE.reg_r17_q , \u_issue.u_regfile.REGFILE.reg_r18_q , \u_issue.u_regfile.REGFILE.reg_r19_q , \u_issue.u_regfile.REGFILE.reg_r20_q , \u_issue.u_regfile.REGFILE.reg_r21_q , \u_issue.u_regfile.REGFILE.reg_r22_q , \u_issue.u_regfile.REGFILE.reg_r23_q , \u_issue.u_regfile.REGFILE.reg_r24_q , \u_issue.u_regfile.REGFILE.reg_r25_q , \u_issue.u_regfile.REGFILE.reg_r26_q , \u_issue.u_regfile.REGFILE.reg_r27_q , \u_issue.u_regfile.REGFILE.reg_r28_q , \u_issue.u_regfile.REGFILE.reg_r29_q , \u_issue.u_regfile.REGFILE.reg_r30_q , \u_issue.u_regfile.REGFILE.reg_r31_q };
  logic [30:0] fangyuan384;
  assign fangyuan384 = { _3815_, _3814_, _3813_, _3812_, _3811_, _3810_, _3809_, _3808_, _3807_, _3806_, _3805_, _3804_, _3803_, _3802_, _3801_, _3800_, _3799_, _3798_, _3797_, _3796_, _3795_, _3794_, _3793_, _3792_, _3791_, _3790_, _3789_, _3788_, _3787_, _3786_, _3785_ };
  always @(32'h00000000 or fangyuan383 or fangyuan384) begin
    casez (fangyuan384)
      31'b??????????????????????????????1 :
        \u_issue.issue_b_rb_value_w = fangyuan383 [31:0] ;
      31'b?????????????????????????????1? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [63:32] ;
      31'b????????????????????????????1?? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [95:64] ;
      31'b???????????????????????????1??? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [127:96] ;
      31'b??????????????????????????1???? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [159:128] ;
      31'b?????????????????????????1????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [191:160] ;
      31'b????????????????????????1?????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [223:192] ;
      31'b???????????????????????1??????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [255:224] ;
      31'b??????????????????????1???????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [287:256] ;
      31'b?????????????????????1????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [319:288] ;
      31'b????????????????????1?????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [351:320] ;
      31'b???????????????????1??????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [383:352] ;
      31'b??????????????????1???????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [415:384] ;
      31'b?????????????????1????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [447:416] ;
      31'b????????????????1?????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [479:448] ;
      31'b???????????????1??????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [511:480] ;
      31'b??????????????1???????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [543:512] ;
      31'b?????????????1????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [575:544] ;
      31'b????????????1?????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [607:576] ;
      31'b???????????1??????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [639:608] ;
      31'b??????????1???????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [671:640] ;
      31'b?????????1????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [703:672] ;
      31'b????????1?????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [735:704] ;
      31'b???????1??????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [767:736] ;
      31'b??????1???????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [799:768] ;
      31'b?????1????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [831:800] ;
      31'b????1?????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [863:832] ;
      31'b???1??????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [895:864] ;
      31'b??1???????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [927:896] ;
      31'b?1????????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [959:928] ;
      31'b1?????????????????????????????? :
        \u_issue.issue_b_rb_value_w = fangyuan383 [991:960] ;
      default:
        \u_issue.issue_b_rb_value_w = 32'h00000000 ;
    endcase
  end
  assign _3785_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1f;
  assign _3786_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1e;
  assign _3787_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1d;
  assign _3788_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1c;
  assign _3789_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1b;
  assign _3790_ = \u_exec1.opcode_opcode_i [24:20] == 5'h1a;
  assign _3791_ = \u_exec1.opcode_opcode_i [24:20] == 5'h19;
  assign _3792_ = \u_exec1.opcode_opcode_i [24:20] == 5'h18;
  assign _3793_ = \u_exec1.opcode_opcode_i [24:20] == 5'h17;
  assign _3794_ = \u_exec1.opcode_opcode_i [24:20] == 5'h16;
  assign _3795_ = \u_exec1.opcode_opcode_i [24:20] == 5'h15;
  assign _3796_ = \u_exec1.opcode_opcode_i [24:20] == 5'h14;
  assign _3797_ = \u_exec1.opcode_opcode_i [24:20] == 5'h13;
  assign _3798_ = \u_exec1.opcode_opcode_i [24:20] == 5'h12;
  assign _3799_ = \u_exec1.opcode_opcode_i [24:20] == 5'h11;
  assign _3800_ = \u_exec1.opcode_opcode_i [24:20] == 5'h10;
  assign _3801_ = \u_exec1.opcode_opcode_i [24:20] == 4'hf;
  assign _3802_ = \u_exec1.opcode_opcode_i [24:20] == 4'he;
  assign _3803_ = \u_exec1.opcode_opcode_i [24:20] == 4'hd;
  assign _3804_ = \u_exec1.opcode_opcode_i [24:20] == 4'hc;
  assign _3805_ = \u_exec1.opcode_opcode_i [24:20] == 4'hb;
  assign _3806_ = \u_exec1.opcode_opcode_i [24:20] == 4'ha;
  assign _3807_ = \u_exec1.opcode_opcode_i [24:20] == 4'h9;
  assign _3808_ = \u_exec1.opcode_opcode_i [24:20] == 4'h8;
  assign _3809_ = \u_exec1.opcode_opcode_i [24:20] == 3'h7;
  assign _3810_ = \u_exec1.opcode_opcode_i [24:20] == 3'h6;
  assign _3811_ = \u_exec1.opcode_opcode_i [24:20] == 3'h5;
  assign _3812_ = \u_exec1.opcode_opcode_i [24:20] == 3'h4;
  assign _3813_ = \u_exec1.opcode_opcode_i [24:20] == 2'h3;
  assign _3814_ = \u_exec1.opcode_opcode_i [24:20] == 2'h2;
  assign _3815_ = \u_exec1.opcode_opcode_i [24:20] == 1'h1;
  logic [991:0] fangyuan385;
  assign fangyuan385 = { \u_issue.u_regfile.REGFILE.reg_r1_q , \u_issue.u_regfile.REGFILE.reg_r2_q , \u_issue.u_regfile.REGFILE.reg_r3_q , \u_issue.u_regfile.REGFILE.reg_r4_q , \u_issue.u_regfile.REGFILE.reg_r5_q , \u_issue.u_regfile.REGFILE.reg_r6_q , \u_issue.u_regfile.REGFILE.reg_r7_q , \u_issue.u_regfile.REGFILE.reg_r8_q , \u_issue.u_regfile.REGFILE.reg_r9_q , \u_issue.u_regfile.REGFILE.reg_r10_q , \u_issue.u_regfile.REGFILE.reg_r11_q , \u_issue.u_regfile.REGFILE.reg_r12_q , \u_issue.u_regfile.REGFILE.reg_r13_q , \u_issue.u_regfile.REGFILE.reg_r14_q , \u_issue.u_regfile.REGFILE.reg_r15_q , \u_issue.u_regfile.REGFILE.reg_r16_q , \u_issue.u_regfile.REGFILE.reg_r17_q , \u_issue.u_regfile.REGFILE.reg_r18_q , \u_issue.u_regfile.REGFILE.reg_r19_q , \u_issue.u_regfile.REGFILE.reg_r20_q , \u_issue.u_regfile.REGFILE.reg_r21_q , \u_issue.u_regfile.REGFILE.reg_r22_q , \u_issue.u_regfile.REGFILE.reg_r23_q , \u_issue.u_regfile.REGFILE.reg_r24_q , \u_issue.u_regfile.REGFILE.reg_r25_q , \u_issue.u_regfile.REGFILE.reg_r26_q , \u_issue.u_regfile.REGFILE.reg_r27_q , \u_issue.u_regfile.REGFILE.reg_r28_q , \u_issue.u_regfile.REGFILE.reg_r29_q , \u_issue.u_regfile.REGFILE.reg_r30_q , \u_issue.u_regfile.REGFILE.reg_r31_q };
  logic [30:0] fangyuan386;
  assign fangyuan386 = { _3846_, _3845_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3838_, _3837_, _3836_, _3835_, _3834_, _3833_, _3832_, _3831_, _3830_, _3829_, _3828_, _3827_, _3826_, _3825_, _3824_, _3823_, _3822_, _3821_, _3820_, _3819_, _3818_, _3817_, _3816_ };
  always @(32'h00000000 or fangyuan385 or fangyuan386) begin
    casez (fangyuan386)
      31'b??????????????????????????????1 :
        \u_issue.issue_b_ra_value_w = fangyuan385 [31:0] ;
      31'b?????????????????????????????1? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [63:32] ;
      31'b????????????????????????????1?? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [95:64] ;
      31'b???????????????????????????1??? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [127:96] ;
      31'b??????????????????????????1???? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [159:128] ;
      31'b?????????????????????????1????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [191:160] ;
      31'b????????????????????????1?????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [223:192] ;
      31'b???????????????????????1??????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [255:224] ;
      31'b??????????????????????1???????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [287:256] ;
      31'b?????????????????????1????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [319:288] ;
      31'b????????????????????1?????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [351:320] ;
      31'b???????????????????1??????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [383:352] ;
      31'b??????????????????1???????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [415:384] ;
      31'b?????????????????1????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [447:416] ;
      31'b????????????????1?????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [479:448] ;
      31'b???????????????1??????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [511:480] ;
      31'b??????????????1???????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [543:512] ;
      31'b?????????????1????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [575:544] ;
      31'b????????????1?????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [607:576] ;
      31'b???????????1??????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [639:608] ;
      31'b??????????1???????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [671:640] ;
      31'b?????????1????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [703:672] ;
      31'b????????1?????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [735:704] ;
      31'b???????1??????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [767:736] ;
      31'b??????1???????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [799:768] ;
      31'b?????1????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [831:800] ;
      31'b????1?????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [863:832] ;
      31'b???1??????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [895:864] ;
      31'b??1???????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [927:896] ;
      31'b?1????????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [959:928] ;
      31'b1?????????????????????????????? :
        \u_issue.issue_b_ra_value_w = fangyuan385 [991:960] ;
      default:
        \u_issue.issue_b_ra_value_w = 32'h00000000 ;
    endcase
  end
  assign _3816_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1f;
  assign _3817_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1e;
  assign _3818_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1d;
  assign _3819_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1c;
  assign _3820_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1b;
  assign _3821_ = \u_exec1.opcode_opcode_i [19:15] == 5'h1a;
  assign _3822_ = \u_exec1.opcode_opcode_i [19:15] == 5'h19;
  assign _3823_ = \u_exec1.opcode_opcode_i [19:15] == 5'h18;
  assign _3824_ = \u_exec1.opcode_opcode_i [19:15] == 5'h17;
  assign _3825_ = \u_exec1.opcode_opcode_i [19:15] == 5'h16;
  assign _3826_ = \u_exec1.opcode_opcode_i [19:15] == 5'h15;
  assign _3827_ = \u_exec1.opcode_opcode_i [19:15] == 5'h14;
  assign _3828_ = \u_exec1.opcode_opcode_i [19:15] == 5'h13;
  assign _3829_ = \u_exec1.opcode_opcode_i [19:15] == 5'h12;
  assign _3830_ = \u_exec1.opcode_opcode_i [19:15] == 5'h11;
  assign _3831_ = \u_exec1.opcode_opcode_i [19:15] == 5'h10;
  assign _3832_ = \u_exec1.opcode_opcode_i [19:15] == 4'hf;
  assign _3833_ = \u_exec1.opcode_opcode_i [19:15] == 4'he;
  assign _3834_ = \u_exec1.opcode_opcode_i [19:15] == 4'hd;
  assign _3835_ = \u_exec1.opcode_opcode_i [19:15] == 4'hc;
  assign _3836_ = \u_exec1.opcode_opcode_i [19:15] == 4'hb;
  assign _3837_ = \u_exec1.opcode_opcode_i [19:15] == 4'ha;
  assign _3838_ = \u_exec1.opcode_opcode_i [19:15] == 4'h9;
  assign _3839_ = \u_exec1.opcode_opcode_i [19:15] == 4'h8;
  assign _3840_ = \u_exec1.opcode_opcode_i [19:15] == 3'h7;
  assign _3841_ = \u_exec1.opcode_opcode_i [19:15] == 3'h6;
  assign _3842_ = \u_exec1.opcode_opcode_i [19:15] == 3'h5;
  assign _3843_ = \u_exec1.opcode_opcode_i [19:15] == 3'h4;
  assign _3844_ = \u_exec1.opcode_opcode_i [19:15] == 2'h3;
  assign _3845_ = \u_exec1.opcode_opcode_i [19:15] == 2'h2;
  assign _3846_ = \u_exec1.opcode_opcode_i [19:15] == 1'h1;
  logic [991:0] fangyuan387;
  assign fangyuan387 = { \u_issue.u_regfile.REGFILE.reg_r1_q , \u_issue.u_regfile.REGFILE.reg_r2_q , \u_issue.u_regfile.REGFILE.reg_r3_q , \u_issue.u_regfile.REGFILE.reg_r4_q , \u_issue.u_regfile.REGFILE.reg_r5_q , \u_issue.u_regfile.REGFILE.reg_r6_q , \u_issue.u_regfile.REGFILE.reg_r7_q , \u_issue.u_regfile.REGFILE.reg_r8_q , \u_issue.u_regfile.REGFILE.reg_r9_q , \u_issue.u_regfile.REGFILE.reg_r10_q , \u_issue.u_regfile.REGFILE.reg_r11_q , \u_issue.u_regfile.REGFILE.reg_r12_q , \u_issue.u_regfile.REGFILE.reg_r13_q , \u_issue.u_regfile.REGFILE.reg_r14_q , \u_issue.u_regfile.REGFILE.reg_r15_q , \u_issue.u_regfile.REGFILE.reg_r16_q , \u_issue.u_regfile.REGFILE.reg_r17_q , \u_issue.u_regfile.REGFILE.reg_r18_q , \u_issue.u_regfile.REGFILE.reg_r19_q , \u_issue.u_regfile.REGFILE.reg_r20_q , \u_issue.u_regfile.REGFILE.reg_r21_q , \u_issue.u_regfile.REGFILE.reg_r22_q , \u_issue.u_regfile.REGFILE.reg_r23_q , \u_issue.u_regfile.REGFILE.reg_r24_q , \u_issue.u_regfile.REGFILE.reg_r25_q , \u_issue.u_regfile.REGFILE.reg_r26_q , \u_issue.u_regfile.REGFILE.reg_r27_q , \u_issue.u_regfile.REGFILE.reg_r28_q , \u_issue.u_regfile.REGFILE.reg_r29_q , \u_issue.u_regfile.REGFILE.reg_r30_q , \u_issue.u_regfile.REGFILE.reg_r31_q };
  logic [30:0] fangyuan388;
  assign fangyuan388 = { _3877_, _3876_, _3875_, _3874_, _3873_, _3872_, _3871_, _3870_, _3869_, _3868_, _3867_, _3866_, _3865_, _3864_, _3863_, _3862_, _3861_, _3860_, _3859_, _3858_, _3857_, _3856_, _3855_, _3854_, _3853_, _3852_, _3851_, _3850_, _3849_, _3848_, _3847_ };
  always @(32'h00000000 or fangyuan387 or fangyuan388) begin
    casez (fangyuan388)
      31'b??????????????????????????????1 :
        \u_issue.issue_a_rb_value_w = fangyuan387 [31:0] ;
      31'b?????????????????????????????1? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [63:32] ;
      31'b????????????????????????????1?? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [95:64] ;
      31'b???????????????????????????1??? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [127:96] ;
      31'b??????????????????????????1???? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [159:128] ;
      31'b?????????????????????????1????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [191:160] ;
      31'b????????????????????????1?????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [223:192] ;
      31'b???????????????????????1??????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [255:224] ;
      31'b??????????????????????1???????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [287:256] ;
      31'b?????????????????????1????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [319:288] ;
      31'b????????????????????1?????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [351:320] ;
      31'b???????????????????1??????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [383:352] ;
      31'b??????????????????1???????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [415:384] ;
      31'b?????????????????1????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [447:416] ;
      31'b????????????????1?????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [479:448] ;
      31'b???????????????1??????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [511:480] ;
      31'b??????????????1???????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [543:512] ;
      31'b?????????????1????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [575:544] ;
      31'b????????????1?????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [607:576] ;
      31'b???????????1??????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [639:608] ;
      31'b??????????1???????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [671:640] ;
      31'b?????????1????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [703:672] ;
      31'b????????1?????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [735:704] ;
      31'b???????1??????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [767:736] ;
      31'b??????1???????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [799:768] ;
      31'b?????1????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [831:800] ;
      31'b????1?????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [863:832] ;
      31'b???1??????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [895:864] ;
      31'b??1???????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [927:896] ;
      31'b?1????????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [959:928] ;
      31'b1?????????????????????????????? :
        \u_issue.issue_a_rb_value_w = fangyuan387 [991:960] ;
      default:
        \u_issue.issue_a_rb_value_w = 32'h00000000 ;
    endcase
  end
  assign _3847_ = \u_csr.opcode_opcode_i [24:20] == 5'h1f;
  assign _3848_ = \u_csr.opcode_opcode_i [24:20] == 5'h1e;
  assign _3849_ = \u_csr.opcode_opcode_i [24:20] == 5'h1d;
  assign _3850_ = \u_csr.opcode_opcode_i [24:20] == 5'h1c;
  assign _3851_ = \u_csr.opcode_opcode_i [24:20] == 5'h1b;
  assign _3852_ = \u_csr.opcode_opcode_i [24:20] == 5'h1a;
  assign _3853_ = \u_csr.opcode_opcode_i [24:20] == 5'h19;
  assign _3854_ = \u_csr.opcode_opcode_i [24:20] == 5'h18;
  assign _3855_ = \u_csr.opcode_opcode_i [24:20] == 5'h17;
  assign _3856_ = \u_csr.opcode_opcode_i [24:20] == 5'h16;
  assign _3857_ = \u_csr.opcode_opcode_i [24:20] == 5'h15;
  assign _3858_ = \u_csr.opcode_opcode_i [24:20] == 5'h14;
  assign _3859_ = \u_csr.opcode_opcode_i [24:20] == 5'h13;
  assign _3860_ = \u_csr.opcode_opcode_i [24:20] == 5'h12;
  assign _3861_ = \u_csr.opcode_opcode_i [24:20] == 5'h11;
  assign _3862_ = \u_csr.opcode_opcode_i [24:20] == 5'h10;
  assign _3863_ = \u_csr.opcode_opcode_i [24:20] == 4'hf;
  assign _3864_ = \u_csr.opcode_opcode_i [24:20] == 4'he;
  assign _3865_ = \u_csr.opcode_opcode_i [24:20] == 4'hd;
  assign _3866_ = \u_csr.opcode_opcode_i [24:20] == 4'hc;
  assign _3867_ = \u_csr.opcode_opcode_i [24:20] == 4'hb;
  assign _3868_ = \u_csr.opcode_opcode_i [24:20] == 4'ha;
  assign _3869_ = \u_csr.opcode_opcode_i [24:20] == 4'h9;
  assign _3870_ = \u_csr.opcode_opcode_i [24:20] == 4'h8;
  assign _3871_ = \u_csr.opcode_opcode_i [24:20] == 3'h7;
  assign _3872_ = \u_csr.opcode_opcode_i [24:20] == 3'h6;
  assign _3873_ = \u_csr.opcode_opcode_i [24:20] == 3'h5;
  assign _3874_ = \u_csr.opcode_opcode_i [24:20] == 3'h4;
  assign _3875_ = \u_csr.opcode_opcode_i [24:20] == 2'h3;
  assign _3876_ = \u_csr.opcode_opcode_i [24:20] == 2'h2;
  assign _3877_ = \u_csr.opcode_opcode_i [24:20] == 1'h1;
  logic [991:0] fangyuan389;
  assign fangyuan389 = { \u_issue.u_regfile.REGFILE.reg_r1_q , \u_issue.u_regfile.REGFILE.reg_r2_q , \u_issue.u_regfile.REGFILE.reg_r3_q , \u_issue.u_regfile.REGFILE.reg_r4_q , \u_issue.u_regfile.REGFILE.reg_r5_q , \u_issue.u_regfile.REGFILE.reg_r6_q , \u_issue.u_regfile.REGFILE.reg_r7_q , \u_issue.u_regfile.REGFILE.reg_r8_q , \u_issue.u_regfile.REGFILE.reg_r9_q , \u_issue.u_regfile.REGFILE.reg_r10_q , \u_issue.u_regfile.REGFILE.reg_r11_q , \u_issue.u_regfile.REGFILE.reg_r12_q , \u_issue.u_regfile.REGFILE.reg_r13_q , \u_issue.u_regfile.REGFILE.reg_r14_q , \u_issue.u_regfile.REGFILE.reg_r15_q , \u_issue.u_regfile.REGFILE.reg_r16_q , \u_issue.u_regfile.REGFILE.reg_r17_q , \u_issue.u_regfile.REGFILE.reg_r18_q , \u_issue.u_regfile.REGFILE.reg_r19_q , \u_issue.u_regfile.REGFILE.reg_r20_q , \u_issue.u_regfile.REGFILE.reg_r21_q , \u_issue.u_regfile.REGFILE.reg_r22_q , \u_issue.u_regfile.REGFILE.reg_r23_q , \u_issue.u_regfile.REGFILE.reg_r24_q , \u_issue.u_regfile.REGFILE.reg_r25_q , \u_issue.u_regfile.REGFILE.reg_r26_q , \u_issue.u_regfile.REGFILE.reg_r27_q , \u_issue.u_regfile.REGFILE.reg_r28_q , \u_issue.u_regfile.REGFILE.reg_r29_q , \u_issue.u_regfile.REGFILE.reg_r30_q , \u_issue.u_regfile.REGFILE.reg_r31_q };
  logic [30:0] fangyuan390;
  assign fangyuan390 = { _3908_, _3907_, _3906_, _3905_, _3904_, _3903_, _3902_, _3901_, _3900_, _3899_, _3898_, _3897_, _3896_, _3895_, _3894_, _3893_, _3892_, _3891_, _3890_, _3889_, _3888_, _3887_, _3886_, _3885_, _3884_, _3883_, _3882_, _3881_, _3880_, _3879_, _3878_ };
  always @(32'h00000000 or fangyuan389 or fangyuan390) begin
    casez (fangyuan390)
      31'b??????????????????????????????1 :
        \u_issue.issue_a_ra_value_w = fangyuan389 [31:0] ;
      31'b?????????????????????????????1? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [63:32] ;
      31'b????????????????????????????1?? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [95:64] ;
      31'b???????????????????????????1??? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [127:96] ;
      31'b??????????????????????????1???? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [159:128] ;
      31'b?????????????????????????1????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [191:160] ;
      31'b????????????????????????1?????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [223:192] ;
      31'b???????????????????????1??????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [255:224] ;
      31'b??????????????????????1???????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [287:256] ;
      31'b?????????????????????1????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [319:288] ;
      31'b????????????????????1?????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [351:320] ;
      31'b???????????????????1??????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [383:352] ;
      31'b??????????????????1???????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [415:384] ;
      31'b?????????????????1????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [447:416] ;
      31'b????????????????1?????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [479:448] ;
      31'b???????????????1??????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [511:480] ;
      31'b??????????????1???????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [543:512] ;
      31'b?????????????1????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [575:544] ;
      31'b????????????1?????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [607:576] ;
      31'b???????????1??????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [639:608] ;
      31'b??????????1???????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [671:640] ;
      31'b?????????1????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [703:672] ;
      31'b????????1?????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [735:704] ;
      31'b???????1??????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [767:736] ;
      31'b??????1???????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [799:768] ;
      31'b?????1????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [831:800] ;
      31'b????1?????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [863:832] ;
      31'b???1??????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [895:864] ;
      31'b??1???????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [927:896] ;
      31'b?1????????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [959:928] ;
      31'b1?????????????????????????????? :
        \u_issue.issue_a_ra_value_w = fangyuan389 [991:960] ;
      default:
        \u_issue.issue_a_ra_value_w = 32'h00000000 ;
    endcase
  end
  assign _3878_ = \u_csr.opcode_opcode_i [19:15] == 5'h1f;
  assign _3879_ = \u_csr.opcode_opcode_i [19:15] == 5'h1e;
  assign _3880_ = \u_csr.opcode_opcode_i [19:15] == 5'h1d;
  assign _3881_ = \u_csr.opcode_opcode_i [19:15] == 5'h1c;
  assign _3882_ = \u_csr.opcode_opcode_i [19:15] == 5'h1b;
  assign _3883_ = \u_csr.opcode_opcode_i [19:15] == 5'h1a;
  assign _3884_ = \u_csr.opcode_opcode_i [19:15] == 5'h19;
  assign _3885_ = \u_csr.opcode_opcode_i [19:15] == 5'h18;
  assign _3886_ = \u_csr.opcode_opcode_i [19:15] == 5'h17;
  assign _3887_ = \u_csr.opcode_opcode_i [19:15] == 5'h16;
  assign _3888_ = \u_csr.opcode_opcode_i [19:15] == 5'h15;
  assign _3889_ = \u_csr.opcode_opcode_i [19:15] == 5'h14;
  assign _3890_ = \u_csr.opcode_opcode_i [19:15] == 5'h13;
  assign _3891_ = \u_csr.opcode_opcode_i [19:15] == 5'h12;
  assign _3892_ = \u_csr.opcode_opcode_i [19:15] == 5'h11;
  assign _3893_ = \u_csr.opcode_opcode_i [19:15] == 5'h10;
  assign _3894_ = \u_csr.opcode_opcode_i [19:15] == 4'hf;
  assign _3895_ = \u_csr.opcode_opcode_i [19:15] == 4'he;
  assign _3896_ = \u_csr.opcode_opcode_i [19:15] == 4'hd;
  assign _3897_ = \u_csr.opcode_opcode_i [19:15] == 4'hc;
  assign _3898_ = \u_csr.opcode_opcode_i [19:15] == 4'hb;
  assign _3899_ = \u_csr.opcode_opcode_i [19:15] == 4'ha;
  assign _3900_ = \u_csr.opcode_opcode_i [19:15] == 4'h9;
  assign _3901_ = \u_csr.opcode_opcode_i [19:15] == 4'h8;
  assign _3902_ = \u_csr.opcode_opcode_i [19:15] == 3'h7;
  assign _3903_ = \u_csr.opcode_opcode_i [19:15] == 3'h6;
  assign _3904_ = \u_csr.opcode_opcode_i [19:15] == 3'h5;
  assign _3905_ = \u_csr.opcode_opcode_i [19:15] == 3'h4;
  assign _3906_ = \u_csr.opcode_opcode_i [19:15] == 2'h3;
  assign _3907_ = \u_csr.opcode_opcode_i [19:15] == 2'h2;
  assign _3908_ = \u_csr.opcode_opcode_i [19:15] == 1'h1;
  assign _3909_ = _3784_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r31_q ;
  assign _3910_ = _3783_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3909_;
  assign _3715_ = rst_i ? 32'h00000000 : _3910_;
  assign _3911_ = _3782_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r30_q ;
  assign _3912_ = _3781_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3911_;
  assign _3714_ = rst_i ? 32'h00000000 : _3912_;
  assign _3913_ = _3780_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r29_q ;
  assign _3914_ = _3779_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3913_;
  assign _3712_ = rst_i ? 32'h00000000 : _3914_;
  assign _3915_ = _3778_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r28_q ;
  assign _3916_ = _3777_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3915_;
  assign _3711_ = rst_i ? 32'h00000000 : _3916_;
  assign _3917_ = _3776_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r27_q ;
  assign _3918_ = _3775_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3917_;
  assign _3710_ = rst_i ? 32'h00000000 : _3918_;
  assign _3919_ = _3774_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r26_q ;
  assign _3920_ = _3773_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3919_;
  assign _3709_ = rst_i ? 32'h00000000 : _3920_;
  assign _3921_ = _3772_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r25_q ;
  assign _3922_ = _3771_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3921_;
  assign _3708_ = rst_i ? 32'h00000000 : _3922_;
  assign _3923_ = _3770_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r24_q ;
  assign _3924_ = _3769_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3923_;
  assign _3707_ = rst_i ? 32'h00000000 : _3924_;
  assign _3925_ = _3768_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r23_q ;
  assign _3926_ = _3767_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3925_;
  assign _3706_ = rst_i ? 32'h00000000 : _3926_;
  assign _3927_ = _3766_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r22_q ;
  assign _3928_ = _3765_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3927_;
  assign _3705_ = rst_i ? 32'h00000000 : _3928_;
  assign _3929_ = _3764_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r21_q ;
  assign _3930_ = _3763_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3929_;
  assign _3704_ = rst_i ? 32'h00000000 : _3930_;
  assign _3931_ = _3762_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r20_q ;
  assign _3932_ = _3761_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3931_;
  assign _3703_ = rst_i ? 32'h00000000 : _3932_;
  assign _3933_ = _3760_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r19_q ;
  assign _3934_ = _3759_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3933_;
  assign _3701_ = rst_i ? 32'h00000000 : _3934_;
  assign _3935_ = _3758_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r18_q ;
  assign _3936_ = _3757_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3935_;
  assign _3700_ = rst_i ? 32'h00000000 : _3936_;
  assign _3937_ = _3756_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r17_q ;
  assign _3938_ = _3755_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3937_;
  assign _3699_ = rst_i ? 32'h00000000 : _3938_;
  assign _3939_ = _3754_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r16_q ;
  assign _3940_ = _3753_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3939_;
  assign _3698_ = rst_i ? 32'h00000000 : _3940_;
  assign _3941_ = _3752_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r15_q ;
  assign _3942_ = _3751_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3941_;
  assign _3697_ = rst_i ? 32'h00000000 : _3942_;
  assign _3943_ = _3750_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r14_q ;
  assign _3944_ = _3749_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3943_;
  assign _3696_ = rst_i ? 32'h00000000 : _3944_;
  assign _3945_ = _3748_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r13_q ;
  assign _3946_ = _3747_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3945_;
  assign _3695_ = rst_i ? 32'h00000000 : _3946_;
  assign _3947_ = _3746_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r12_q ;
  assign _3948_ = _3745_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3947_;
  assign _3694_ = rst_i ? 32'h00000000 : _3948_;
  assign _3949_ = _3744_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r11_q ;
  assign _3950_ = _3743_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3949_;
  assign _3693_ = rst_i ? 32'h00000000 : _3950_;
  assign _3951_ = _3742_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r10_q ;
  assign _3952_ = _3741_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3951_;
  assign _3692_ = rst_i ? 32'h00000000 : _3952_;
  assign _3953_ = _3740_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r9_q ;
  assign _3954_ = _3739_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3953_;
  assign _3722_ = rst_i ? 32'h00000000 : _3954_;
  assign _3955_ = _3738_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r8_q ;
  assign _3956_ = _3737_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3955_;
  assign _3721_ = rst_i ? 32'h00000000 : _3956_;
  assign _3957_ = _3736_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r7_q ;
  assign _3958_ = _3735_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3957_;
  assign _3720_ = rst_i ? 32'h00000000 : _3958_;
  assign _3959_ = _3734_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r6_q ;
  assign _3960_ = _3733_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3959_;
  assign _3719_ = rst_i ? 32'h00000000 : _3960_;
  assign _3961_ = _3732_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r5_q ;
  assign _3962_ = _3731_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3961_;
  assign _3718_ = rst_i ? 32'h00000000 : _3962_;
  assign _3963_ = _3730_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r4_q ;
  assign _3964_ = _3729_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3963_;
  assign _3717_ = rst_i ? 32'h00000000 : _3964_;
  assign _3965_ = _3728_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r3_q ;
  assign _3966_ = _3727_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3965_;
  assign _3716_ = rst_i ? 32'h00000000 : _3966_;
  assign _3967_ = _3726_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r2_q ;
  assign _3968_ = _3725_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3967_;
  assign _3713_ = rst_i ? 32'h00000000 : _3968_;
  assign _3969_ = _3724_ ? \u_issue.u_pipe1_ctrl.result_wb_q : \u_issue.u_regfile.REGFILE.reg_r1_q ;
  assign _3970_ = _3723_ ? \u_issue.u_pipe0_ctrl.result_wb_q : _3969_;
  assign _3702_ = rst_i ? 32'h00000000 : _3970_;
  logic [31:0] fangyuan391;
  assign fangyuan391 = { \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31:20] };
  assign _4003_ = \u_issue.lsu_opcode_ra_operand_o + fangyuan391;
  logic [31:0] fangyuan392;
  assign fangyuan392 = { \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31], \u_issue.lsu_opcode_opcode_o [31:25], \u_issue.lsu_opcode_opcode_o [11:7] };
  assign _4004_ = \u_issue.lsu_opcode_ra_operand_o + fangyuan392;
  assign \u_lsu.complete_ok_e2_w = mem_d_ack_i & _4071_;
  assign \u_lsu.complete_err_e2_w = mem_d_ack_i & mem_d_error_i;
  assign _4005_ = \u_lsu.mem_unaligned_e1_q & _4072_;
  assign _4006_ = \u_issue.lsu_opcode_opcode_o & 15'h707f;
  assign _4007_ = \u_issue.lsu_opcode_valid_o & \u_lsu.dcache_invalidate_w ;
  assign _4008_ = \u_issue.lsu_opcode_valid_o & \u_lsu.dcache_writeback_w ;
  assign _4009_ = \u_issue.lsu_opcode_valid_o & \u_lsu.dcache_flush_w ;
  assign \u_lsu.mem_rd_o = \u_lsu.mem_rd_q & _4072_;
  assign \u_lsu.mem_wr_o = \u_lsu.mem_wr_q & _4073_;
  assign \u_lsu.fault_load_align_w = \u_lsu.mem_unaligned_e2_q & \u_lsu.u_lsu_request.data_out_o [0];
  assign \u_lsu.fault_store_align_w = \u_lsu.mem_unaligned_e2_q & _4074_;
  assign _4013_ = _4006_ == 2'h3;
  assign _4014_ = _4006_ == 13'h1003;
  assign _4015_ = _4006_ == 14'h2003;
  assign _4016_ = _4006_ == 15'h4003;
  assign _4017_ = _4006_ == 15'h5003;
  assign _4018_ = _4006_ == 15'h6003;
  assign \u_lsu.req_sb_w = _4006_ == 6'h23;
  assign \u_lsu.req_sh_w = _4006_ == 13'h1023;
  assign _4019_ = _4006_ == 14'h2023;
  assign _4020_ = _4006_ == 13'h1073;
  assign _4021_ = \u_issue.lsu_opcode_opcode_o [31:20] == 10'h3a0;
  assign _4022_ = \u_issue.lsu_opcode_opcode_o [31:20] == 10'h3a1;
  assign _4023_ = \u_issue.lsu_opcode_opcode_o [31:20] == 10'h3a2;
  assign _4024_ = \u_lsu.mem_addr_r >= 32'h80000000;
  assign _4025_ = \u_lsu.mem_addr_r <= 32'h8fffffff;
  assign \u_lsu.issue_lsu_e1_w = _4050_ && mem_d_accept_i;
  assign \u_lsu.delay_lsu_e2_w = \u_lsu.pending_lsu_e2_q && _4044_;
  assign _4026_ = \u_issue.lsu_opcode_valid_o && _4020_;
  assign _4027_ = \u_issue.lsu_opcode_valid_o && \u_lsu.load_inst_w ;
  assign _4028_ = \u_issue.lsu_opcode_valid_o && \u_lsu.req_sw_lw_w ;
  assign _4029_ = \u_issue.lsu_opcode_valid_o && \u_lsu.req_sh_lh_w ;
  assign \u_lsu.mem_rd_r = _4027_ && _4045_;
  assign _4030_ = \u_issue.lsu_opcode_valid_o && _4019_;
  assign _4031_ = _4030_ && _4045_;
  assign _4032_ = \u_issue.lsu_opcode_valid_o && \u_lsu.req_sh_w ;
  assign _4033_ = _4032_ && _4045_;
  assign _4034_ = \u_issue.lsu_opcode_valid_o && \u_lsu.req_sb_w ;
  assign \u_lsu.dcache_flush_w = _4020_ && _4021_;
  assign \u_lsu.dcache_writeback_w = _4020_ && _4022_;
  assign \u_lsu.dcache_invalidate_w = _4020_ && _4023_;
  assign _4035_ = _4059_ && \u_lsu.delay_lsu_e2_w ;
  assign _4036_ = _4063_ && _4046_;
  assign _4037_ = _4024_ && _4025_;
  assign _4038_ = \u_issue.lsu_opcode_valid_o && _4065_;
  assign _4039_ = \u_lsu.mem_unaligned_e1_q && _4072_;
  assign _4040_ = mem_d_ack_i && mem_d_error_i;
  assign _4041_ = mem_d_ack_i && \u_lsu.u_lsu_request.data_out_o [0];
  assign _4042_ = \u_lsu.u_lsu_request.data_out_o [3] && _3996_[7];
  assign _4043_ = \u_lsu.u_lsu_request.data_out_o [3] && _4001_[15];
  assign \u_lsu.fault_load_bus_w = mem_d_error_i && \u_lsu.u_lsu_request.data_out_o [0];
  assign \u_lsu.fault_store_bus_w = mem_d_error_i && _4074_;
  assign \u_lsu.fault_load_page_w = mem_d_error_i && 1'h0;
  assign \u_lsu.fault_store_page_w = mem_d_error_i && 1'h0;
  assign _4044_ = ! \u_lsu.complete_ok_e2_w ;
  assign _4045_ = ! \u_lsu.mem_unaligned_r ;
  assign _4046_ = ! mem_d_accept_i;
  assign _4047_ = \u_lsu.mem_rd_o || _4126_;
  assign _4048_ = _4047_ || \u_lsu.mem_writeback_q ;
  assign _4049_ = _4048_ || \u_lsu.mem_invalidate_q ;
  assign _4050_ = _4049_ || \u_lsu.mem_flush_q ;
  assign _4051_ = \u_lsu.complete_ok_e2_w || \u_lsu.complete_err_e2_w ;
  assign _4052_ = _4013_ || _4014_;
  assign \u_lsu.load_signed_inst_w = _4052_ || _4015_;
  assign _4053_ = \u_lsu.load_signed_inst_w || _4016_;
  assign _4054_ = _4053_ || _4017_;
  assign \u_lsu.load_inst_w = _4054_ || _4018_;
  assign \u_lsu.req_lb_w = _4013_ || _4016_;
  assign \u_lsu.req_lh_w = _4014_ || _4017_;
  assign _4055_ = _4019_ || _4015_;
  assign \u_lsu.req_sw_lw_w = _4055_ || _4018_;
  assign _4056_ = \u_lsu.req_sh_w || _4014_;
  assign \u_lsu.req_sh_lh_w = _4056_ || _4017_;
  assign _4057_ = \u_lsu.complete_err_e2_w || \u_lsu.mem_unaligned_e2_q ;
  assign _4058_ = \u_lsu.mem_rd_q || _4127_;
  assign _4059_ = _4058_ || \u_lsu.mem_unaligned_e1_q ;
  assign _4060_ = \u_lsu.mem_writeback_q || \u_lsu.mem_invalidate_q ;
  assign _4061_ = _4060_ || \u_lsu.mem_flush_q ;
  assign _4062_ = _4061_ || \u_lsu.mem_rd_o ;
  assign _4063_ = _4062_ || _4070_;
  assign _4064_ = \u_lsu.dcache_invalidate_w || \u_lsu.dcache_writeback_w ;
  assign _4065_ = _4064_ || \u_lsu.dcache_flush_w ;
  assign _4066_ = _4037_ || _4038_;
  assign _4067_ = _4036_ || \u_lsu.delay_lsu_e2_w ;
  assign \u_issue.lsu_stall_i = _4067_ || \u_lsu.mem_unaligned_e1_q ;
  assign \u_lsu.u_lsu_request.push_i = \u_lsu.issue_lsu_e1_w || _4039_;
  assign \u_lsu.u_lsu_request.pop_i = mem_d_ack_i || \u_lsu.mem_unaligned_e2_q ;
  assign _4068_ = _4040_ || \u_lsu.mem_unaligned_e2_q ;
  assign _4069_ = | \u_lsu.mem_addr_r [1:0];
  assign _4070_ = | \u_lsu.mem_wr_o ;
  assign _4071_ = ~ mem_d_error_i;
  assign _4072_ = ~ \u_lsu.delay_lsu_e2_w ;
  logic [3:0] fangyuan393;
  assign fangyuan393 = { \u_lsu.delay_lsu_e2_w , \u_lsu.delay_lsu_e2_w , \u_lsu.delay_lsu_e2_w , \u_lsu.delay_lsu_e2_w };
  assign _4073_ = ~ fangyuan393;
  assign _4074_ = ~ \u_lsu.u_lsu_request.data_out_o [0];
  assign _4075_ = \u_lsu.req_lb_w | \u_lsu.req_sb_w ;
  assign _4076_ = \u_lsu.req_lh_w | \u_lsu.req_sh_w ;
  assign \u_issue.u_pipe0_ctrl.mem_complete_i = mem_d_ack_i | \u_lsu.mem_unaligned_e2_q ;
  always @(posedge clk_i)
      \u_lsu.mem_addr_q <= _3971_;
  always @(posedge clk_i)
      \u_lsu.mem_data_wr_q <= _3973_;
  always @(posedge clk_i)
      \u_lsu.mem_rd_q <= _3978_;
  always @(posedge clk_i)
      \u_lsu.mem_wr_q <= _3981_;
  always @(posedge clk_i)
      \u_lsu.mem_cacheable_q <= _3972_;
  always @(posedge clk_i)
      \u_lsu.mem_invalidate_q <= _3975_;
  always @(posedge clk_i)
      \u_lsu.mem_writeback_q <= _3982_;
  always @(posedge clk_i)
      \u_lsu.mem_flush_q <= _3974_;
  always @(posedge clk_i)
      \u_lsu.mem_unaligned_e1_q <= _3979_;
  always @(posedge clk_i)
      \u_lsu.mem_load_q <= _3976_;
  always @(posedge clk_i)
      \u_lsu.mem_xb_q <= _3983_;
  always @(posedge clk_i)
      \u_lsu.mem_xh_q <= _3984_;
  always @(posedge clk_i)
      \u_lsu.mem_ls_q <= _3977_;
  always @(posedge clk_i)
      \u_lsu.mem_unaligned_e2_q <= _3980_;
  always @(posedge clk_i)
      \u_lsu.pending_lsu_e2_q <= _3985_;
  logic [31:0] fangyuan394;
  assign fangyuan394 = { 16'hffff, _4001_ };
  logic [31:0] fangyuan395;
  assign fangyuan395 = { 16'h0000, _4001_ };
  assign _4002_ = _4043_ ? fangyuan394 : fangyuan395;
  assign _4001_ = \u_lsu.u_lsu_request.data_out_o [5] ? mem_d_data_rd_i[31:16] : mem_d_data_rd_i[15:0];
  assign _4000_ = \u_lsu.u_lsu_request.data_out_o [2] ? _4002_ : mem_d_data_rd_i;
  logic [31:0] fangyuan396;
  assign fangyuan396 = { 24'hffffff, _3996_ };
  logic [31:0] fangyuan397;
  assign fangyuan397 = { 24'h000000, _3996_ };
  assign _3999_ = _4042_ ? fangyuan396 : fangyuan397;
  logic [3:0] fangyuan398;
  assign fangyuan398 = { _4080_, _4079_, _4078_, _4077_ };
  always @(8'hxx or mem_d_data_rd_i or fangyuan398) begin
    casez (fangyuan398)
      4'b???1 :
        _3996_ = mem_d_data_rd_i [7:0] ;
      4'b??1? :
        _3996_ = mem_d_data_rd_i [15:8] ;
      4'b?1?? :
        _3996_ = mem_d_data_rd_i [23:16] ;
      4'b1??? :
        _3996_ = mem_d_data_rd_i [31:24] ;
      default:
        _3996_ = 8'hxx ;
    endcase
  end
  assign _4077_ = ! \u_lsu.u_lsu_request.data_out_o [5:4];
  assign _4078_ = \u_lsu.u_lsu_request.data_out_o [5:4] == 1'h1;
  assign _4079_ = \u_lsu.u_lsu_request.data_out_o [5:4] == 2'h2;
  assign _4080_ = \u_lsu.u_lsu_request.data_out_o [5:4] == 2'h3;
  assign _3993_ = \u_lsu.u_lsu_request.data_out_o [1] ? _3999_ : _4000_;
  assign _3990_ = _4041_ ? _3993_ : 32'h00000000;
  assign \u_issue.u_pipe0_ctrl.mem_result_e2_i = _4068_ ? \u_lsu.u_lsu_request.data_out_o [35:4] : _3990_;
  assign _4081_ = _4036_ ? \u_lsu.mem_ls_q : \u_lsu.load_signed_inst_w ;
  assign _4082_ = _4035_ ? \u_lsu.mem_ls_q : _4081_;
  assign _4083_ = _4057_ ? 1'h0 : _4082_;
  assign _3977_ = rst_i ? 1'h0 : _4083_;
  assign _4084_ = _4036_ ? \u_lsu.mem_xh_q : _4076_;
  assign _4085_ = _4035_ ? \u_lsu.mem_xh_q : _4084_;
  assign _4086_ = _4057_ ? 1'h0 : _4085_;
  assign _3984_ = rst_i ? 1'h0 : _4086_;
  assign _4087_ = _4036_ ? \u_lsu.mem_xb_q : _4075_;
  assign _4088_ = _4035_ ? \u_lsu.mem_xb_q : _4087_;
  assign _4089_ = _4057_ ? 1'h0 : _4088_;
  assign _3983_ = rst_i ? 1'h0 : _4089_;
  assign _4090_ = _4036_ ? \u_lsu.mem_load_q : _4027_;
  assign _4091_ = _4035_ ? \u_lsu.mem_load_q : _4090_;
  assign _4092_ = _4057_ ? 1'h0 : _4091_;
  assign _3976_ = rst_i ? 1'h0 : _4092_;
  assign _4093_ = _4036_ ? \u_lsu.mem_unaligned_e1_q : \u_lsu.mem_unaligned_r ;
  assign _4094_ = _4035_ ? \u_lsu.mem_unaligned_e1_q : _4093_;
  assign _4095_ = _4057_ ? 1'h0 : _4094_;
  assign _3979_ = rst_i ? 1'h0 : _4095_;
  assign _4096_ = _4036_ ? \u_lsu.mem_flush_q : _4009_;
  assign _4097_ = _4035_ ? \u_lsu.mem_flush_q : _4096_;
  assign _4098_ = _4057_ ? 1'h0 : _4097_;
  assign _3974_ = rst_i ? 1'h0 : _4098_;
  assign _4099_ = _4036_ ? \u_lsu.mem_writeback_q : _4008_;
  assign _4100_ = _4035_ ? \u_lsu.mem_writeback_q : _4099_;
  assign _4101_ = _4057_ ? 1'h0 : _4100_;
  assign _3982_ = rst_i ? 1'h0 : _4101_;
  assign _4102_ = _4036_ ? \u_lsu.mem_invalidate_q : _4007_;
  assign _4103_ = _4035_ ? \u_lsu.mem_invalidate_q : _4102_;
  assign _4104_ = _4057_ ? 1'h0 : _4103_;
  assign _3975_ = rst_i ? 1'h0 : _4104_;
  assign _4105_ = _4036_ ? \u_lsu.mem_cacheable_q : _4066_;
  assign _4106_ = _4035_ ? \u_lsu.mem_cacheable_q : _4105_;
  assign _4107_ = _4057_ ? 1'h0 : _4106_;
  assign _3972_ = rst_i ? 1'h0 : _4107_;
  assign _4108_ = _4036_ ? \u_lsu.mem_wr_q : \u_lsu.mem_wr_r ;
  assign _4109_ = _4035_ ? \u_lsu.mem_wr_q : _4108_;
  assign _4110_ = _4057_ ? 4'h0 : _4109_;
  assign _3981_ = rst_i ? 4'h0 : _4110_;
  assign _4111_ = _4036_ ? \u_lsu.mem_rd_q : \u_lsu.mem_rd_r ;
  assign _4112_ = _4035_ ? \u_lsu.mem_rd_q : _4111_;
  assign _4113_ = _4057_ ? 1'h0 : _4112_;
  assign _3978_ = rst_i ? 1'h0 : _4113_;
  assign _4114_ = _4036_ ? \u_lsu.mem_data_wr_q : \u_lsu.mem_data_r ;
  assign _4115_ = _4035_ ? \u_lsu.mem_data_wr_q : _4114_;
  assign _4116_ = _4057_ ? 32'h00000000 : _4115_;
  assign _3973_ = rst_i ? 32'h00000000 : _4116_;
  assign _4117_ = _4036_ ? \u_lsu.mem_addr_q : \u_lsu.mem_addr_r ;
  assign _4118_ = _4035_ ? \u_lsu.mem_addr_q : _4117_;
  assign _4119_ = _4057_ ? 32'h00000000 : _4118_;
  assign _3971_ = rst_i ? 32'h00000000 : _4119_;
  logic [3:0] fangyuan399;
  assign fangyuan399 = { _4123_, _4122_, _4121_, _4120_ };
  always @(4'hx or fangyuan399) begin
    casez (fangyuan399)
      4'b???1 :
        _3998_ = 4'b0001 ;
      4'b??1? :
        _3998_ = 4'b0010 ;
      4'b?1?? :
        _3998_ = 4'b0100 ;
      4'b1??? :
        _3998_ = 4'b1000 ;
      default:
        _3998_ = 4'hx ;
    endcase
  end
  assign _4120_ = ! \u_lsu.mem_addr_r [1:0];
  assign _4121_ = \u_lsu.mem_addr_r [1:0] == 1'h1;
  assign _4122_ = \u_lsu.mem_addr_r [1:0] == 2'h2;
  assign _4123_ = \u_lsu.mem_addr_r [1:0] == 2'h3;
  logic [127:0] fangyuan400;
  assign fangyuan400 = { \u_issue.lsu_opcode_rb_operand_o [7:0], 16'h0000, 16'h0000, \u_issue.lsu_opcode_rb_operand_o [7:0], 16'h0000, 16'h0000, \u_issue.lsu_opcode_rb_operand_o [7:0], 16'h0000, 16'h0000, \u_issue.lsu_opcode_rb_operand_o [7:0] };
  logic [3:0] fangyuan401;
  assign fangyuan401 = { _4123_, _4122_, _4121_, _4120_ };
  always @(32'hxxxxxxxx or fangyuan400 or fangyuan401) begin
    casez (fangyuan401)
      4'b???1 :
        _3997_ = fangyuan400 [31:0] ;
      4'b??1? :
        _3997_ = fangyuan400 [63:32] ;
      4'b?1?? :
        _3997_ = fangyuan400 [95:64] ;
      4'b1??? :
        _3997_ = fangyuan400 [127:96] ;
      default:
        _3997_ = 32'hxxxxxxxx ;
    endcase
  end
  assign _3995_ = _4034_ ? _3998_ : 4'h0;
  assign _3994_ = _4034_ ? _3997_ : 32'h00000000;
  assign _3992_ = _4122_ ? 4'hc : 4'h3;
  logic [31:0] fangyuan402;
  assign fangyuan402 = { \u_issue.lsu_opcode_rb_operand_o [15:0], 16'h0000 };
  logic [31:0] fangyuan403;
  assign fangyuan403 = { 16'h0000, \u_issue.lsu_opcode_rb_operand_o [15:0] };
  assign _3991_ = _4122_ ? fangyuan402 : fangyuan403;
  assign _3989_ = _4033_ ? _3992_ : _3995_;
  assign _3987_ = _4033_ ? _3991_ : _3994_;
  assign \u_lsu.mem_wr_r = _4031_ ? 4'hf : _3989_;
  assign \u_lsu.mem_data_r = _4031_ ? \u_issue.lsu_opcode_rb_operand_o : _3987_;
  assign _3988_ = _4029_ ? \u_lsu.mem_addr_r [0] : 1'h0;
  assign \u_lsu.mem_unaligned_r = _4028_ ? _4069_ : _3988_;
  assign _3986_ = _4027_ ? _4003_ : _4004_;
  assign \u_lsu.mem_addr_r = _4026_ ? \u_issue.lsu_opcode_ra_operand_o : _3986_;
  assign _3980_ = rst_i ? 1'h0 : _4005_;
  assign _4124_ = _4051_ ? 1'h0 : \u_lsu.pending_lsu_e2_q ;
  assign _4125_ = \u_lsu.issue_lsu_e1_w ? 1'h1 : _4124_;
  assign _3985_ = rst_i ? 1'h0 : _4125_;
  logic [3:0] fangyuan404;
  assign fangyuan404 = { \u_lsu.mem_wr_o [0], \u_lsu.mem_wr_o [1], \u_lsu.mem_wr_o [2], \u_lsu.mem_wr_o [3] };
  assign _4126_ = | fangyuan404;
  logic [3:0] fangyuan405;
  assign fangyuan405 = { \u_lsu.mem_wr_q [0], \u_lsu.mem_wr_q [1], \u_lsu.mem_wr_q [2], \u_lsu.mem_wr_q [3] };
  assign _4127_ = | fangyuan405;
  assign _4010_[4:0] = \u_lsu.fault_store_bus_w ? 5'h17 : 5'h00;
  assign _4011_[4:0] = \u_lsu.fault_load_bus_w ? 5'h15 : _4010_[4:0];
  assign _4128_[4:0] = \u_lsu.fault_store_page_w ? 5'h1f : _4011_[4:0];
  assign _4012_[4:0] = \u_lsu.fault_load_page_w ? 5'h1d : _4128_[4:0];
  assign _4129_[4:0] = \u_lsu.fault_store_align_w ? 5'h16 : _4012_[4:0];
  assign \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] = \u_lsu.fault_load_align_w ? 5'h14 : _4129_[4:0];
  assign _4135_ = \u_lsu.u_lsu_request.wr_ptr_q + 1'h1;
  assign _4136_[0] = \u_lsu.u_lsu_request.rd_ptr_q + 1'h1;
  assign _4137_ = \u_lsu.u_lsu_request.count_q + 1'h1;
  assign _4138_ = \u_lsu.u_lsu_request.push_i & \u_lsu.u_lsu_request.accept_o ;
  assign _4139_ = \u_lsu.u_lsu_request.pop_i & \u_lsu.u_lsu_request.valid_o ;
  assign _4140_ = _4138_ & _4142_;
  assign _4141_ = _4143_ & _4139_;
  assign \u_lsu.u_lsu_request.valid_o = | \u_lsu.u_lsu_request.count_q ;
  assign \u_lsu.u_lsu_request.accept_o = \u_lsu.u_lsu_request.count_q != 2'h2;
  assign _4142_ = ~ _4139_;
  assign _4143_ = ~ _4138_;
  always @(posedge clk_i)
      \u_lsu.u_lsu_request.rd_ptr_q <= _4133_;
  always @(posedge clk_i)
      \u_lsu.u_lsu_request.wr_ptr_q <= _4134_;
  always @(posedge clk_i)
      \u_lsu.u_lsu_request.count_q <= _4132_;
  assign _4130_[35] = rst_i ? 1'h1 : 1'h0;
  assign _4144_[35] = _4138_ ? 1'h1 : 1'h0;
  assign _4131_[35] = rst_i ? 1'h0 : _4144_[35];
  assign _4145_ = _4141_ ? _4149_[1:0] : \u_lsu.u_lsu_request.count_q ;
  assign _4146_ = _4140_ ? _4137_ : _4145_;
  assign _4132_ = rst_i ? 2'h0 : _4146_;
  assign _4147_ = _4138_ ? _4135_ : \u_lsu.u_lsu_request.wr_ptr_q ;
  assign _4134_ = rst_i ? 1'h0 : _4147_;
  assign _4148_ = _4139_ ? _4136_[0] : \u_lsu.u_lsu_request.rd_ptr_q ;
  assign _4133_ = rst_i ? 1'h0 : _4148_;
  assign _4149_[1:0] = \u_lsu.u_lsu_request.count_q - 1'h1;
  assign _4156_ = \u_issue.mul_opcode_opcode_o & 32'hfe00707f;
  assign _4157_ = _4156_ == 26'h2000033;
  assign _4158_ = _4156_ == 26'h2001033;
  assign _4159_ = _4156_ == 26'h2002033;
  assign _4160_ = _4156_ == 26'h2003033;
  assign _4161_ = \u_issue.mul_opcode_valid_o && \u_mul.mult_inst_w ;
  assign _4162_ = _4157_ || _4158_;
  assign _4163_ = _4162_ || _4159_;
  assign \u_mul.mult_inst_w = _4163_ || _4160_;
  logic [64:0] fangyuan406;
  assign fangyuan406 = { \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q [32], \u_mul.operand_a_e1_q };
  logic [64:0] fangyuan407;
  assign fangyuan407 = { \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q [32], \u_mul.operand_b_e1_q };
  assign \u_mul.mult_result_w = fangyuan406 * fangyuan407;
  assign _4164_ = ~ _4157_;
  always @(posedge clk_i)
      \u_mul.result_e2_q <= _4153_;
  always @(posedge clk_i)
      \u_mul.operand_a_e1_q <= _4151_;
  always @(posedge clk_i)
      \u_mul.operand_b_e1_q <= _4152_;
  always @(posedge clk_i)
      \u_mul.mulhi_sel_e1_q <= _4150_;
  assign _4165_ = \u_exec0.hold_i ? \u_mul.result_e2_q : \u_mul.result_r ;
  assign _4153_ = rst_i ? 32'h00000000 : _4165_;
  assign _4166_ = _4161_ ? _4164_ : 1'h0;
  assign _4167_ = \u_exec0.hold_i ? \u_mul.mulhi_sel_e1_q : _4166_;
  assign _4150_ = rst_i ? 1'h0 : _4167_;
  assign _4168_ = _4161_ ? \u_mul.operand_b_r : 33'h000000000;
  assign _4169_ = \u_exec0.hold_i ? \u_mul.operand_b_e1_q : _4168_;
  assign _4152_ = rst_i ? 33'h000000000 : _4169_;
  assign _4170_ = _4161_ ? \u_mul.operand_a_r : 33'h000000000;
  assign _4171_ = \u_exec0.hold_i ? \u_mul.operand_a_e1_q : _4170_;
  assign _4151_ = rst_i ? 33'h000000000 : _4171_;
  logic [32:0] fangyuan408;
  assign fangyuan408 = { \u_issue.mul_opcode_rb_operand_o [31], \u_issue.mul_opcode_rb_operand_o };
  logic [32:0] fangyuan409;
  assign fangyuan409 = { 1'h0, \u_issue.mul_opcode_rb_operand_o };
  assign _4155_ = _4158_ ? fangyuan408 : fangyuan409;
  logic [32:0] fangyuan410;
  assign fangyuan410 = { 1'h0, \u_issue.mul_opcode_rb_operand_o };
  assign \u_mul.operand_b_r = _4159_ ? fangyuan410 : _4155_;
  logic [32:0] fangyuan411;
  assign fangyuan411 = { \u_issue.mul_opcode_ra_operand_o [31], \u_issue.mul_opcode_ra_operand_o };
  logic [32:0] fangyuan412;
  assign fangyuan412 = { 1'h0, \u_issue.mul_opcode_ra_operand_o };
  assign _4154_ = _4158_ ? fangyuan411 : fangyuan412;
  logic [32:0] fangyuan413;
  assign fangyuan413 = { \u_issue.mul_opcode_ra_operand_o [31], \u_issue.mul_opcode_ra_operand_o };
  assign \u_mul.operand_a_r = _4159_ ? fangyuan413 : _4154_;
  assign \u_mul.result_r = \u_mul.mulhi_sel_e1_q ? \u_mul.mult_result_w [63:32] : \u_mul.mult_result_w [31:0];
  assign branch_csr_pc_w = \u_csr.branch_target_q ;
  assign branch_csr_request_w = \u_csr.branch_q ;
  assign branch_d_exec0_pc_w = \u_exec0.branch_target_r ;
  assign branch_d_exec0_request_w = \u_exec0.branch_d_request_o ;
  assign branch_d_exec1_pc_w = \u_exec1.branch_target_r ;
  assign branch_d_exec1_request_w = \u_exec1.branch_d_request_o ;
  assign branch_exec0_is_call_w = \u_exec0.branch_call_q ;
  assign branch_exec0_is_jmp_w = \u_exec0.branch_jmp_q ;
  assign branch_exec0_is_not_taken_w = \u_exec0.branch_ntaken_q ;
  assign branch_exec0_is_ret_w = \u_exec0.branch_ret_q ;
  assign branch_exec0_is_taken_w = \u_exec0.branch_taken_q ;
  assign branch_exec0_pc_w = \u_exec0.pc_x_q ;
  assign branch_exec0_source_w = \u_exec0.pc_m_q ;
  assign branch_exec1_is_call_w = \u_exec1.branch_call_q ;
  assign branch_exec1_is_jmp_w = \u_exec1.branch_jmp_q ;
  assign branch_exec1_is_not_taken_w = \u_exec1.branch_ntaken_q ;
  assign branch_exec1_is_ret_w = \u_exec1.branch_ret_q ;
  assign branch_exec1_is_taken_w = \u_exec1.branch_taken_q ;
  assign branch_exec1_pc_w = \u_exec1.pc_x_q ;
  assign branch_exec1_request_w = \u_exec1.branch_request_o ;
  assign branch_exec1_source_w = \u_exec1.pc_m_q ;
  assign branch_info_is_call_w = \u_frontend.u_npc.branch_is_call_i ;
  assign branch_info_is_jmp_w = \u_frontend.u_npc.branch_is_jmp_i ;
  assign branch_info_is_not_taken_w = \u_frontend.u_npc.branch_is_not_taken_i ;
  assign branch_info_is_ret_w = \u_frontend.u_npc.branch_is_ret_i ;
  assign branch_info_is_taken_w = \u_frontend.u_npc.branch_is_taken_i ;
  assign branch_info_pc_w = \u_frontend.u_npc.branch_pc_i ;
  assign branch_info_request_w = \u_frontend.u_npc.branch_request_i ;
  assign branch_info_source_w = \u_frontend.u_npc.branch_source_i ;
  assign branch_pc_w = \u_frontend.u_fetch.branch_pc_i ;
  assign branch_request_w = \u_frontend.u_decode.u_fifo.flush_i ;
  assign csr_opcode_invalid_w = \u_csr.opcode_invalid_i ;
  assign csr_opcode_opcode_w = \u_csr.opcode_opcode_i ;
  assign csr_opcode_pc_w = \u_exec0.opcode_pc_i ;
  assign csr_opcode_ra_idx_w = \u_csr.opcode_opcode_i [19:15];
  assign csr_opcode_ra_operand_w = \u_csr.opcode_ra_operand_i ;
  assign csr_opcode_rb_idx_w = \u_csr.opcode_opcode_i [24:20];
  assign csr_opcode_rb_operand_w = \u_div.opcode_rb_operand_i ;
  assign csr_opcode_rd_idx_w = \u_csr.opcode_opcode_i [11:7];
  assign csr_opcode_valid_w = \u_csr.opcode_valid_i ;
  assign csr_result_e1_exception_w = \u_csr.exception_e1_q ;
  assign csr_result_e1_value_w = \u_csr.rd_result_e1_q ;
  assign csr_result_e1_wdata_w = \u_csr.csr_wdata_e1_q ;
  assign csr_result_e1_write_w = \u_csr.rd_valid_e1_q ;
  assign csr_writeback_exception_addr_w = \u_csr.u_csrfile.exception_addr_i ;
  assign csr_writeback_exception_pc_w = \u_csr.u_csrfile.exception_pc_i ;
  assign csr_writeback_exception_w = \u_csr.u_csrfile.exception_i ;
  assign csr_writeback_waddr_w = \u_issue.u_pipe0_ctrl.opcode_wb_q [31:20];
  assign csr_writeback_wdata_w = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  assign csr_writeback_write_w = \u_issue.u_pipe0_ctrl.csr_wr_wb_q ;
  assign div_opcode_valid_w = \u_div.opcode_valid_i ;
  assign exec0_hold_w = \u_exec0.hold_i ;
  assign exec0_opcode_valid_w = \u_div.opcode_valid_i ;
  assign exec1_hold_w = \u_exec0.hold_i ;
  assign exec1_opcode_valid_w = \u_exec1.opcode_valid_i ;
  assign fetch0_accept_w = \u_frontend.u_decode.u_fifo.pop0_i ;
  assign fetch0_fault_fetch_w = \u_frontend.u_decode.u_fifo.info0_out_o [0];
  assign fetch0_fault_page_w = \u_frontend.u_decode.u_fifo.info0_out_o [1];
  assign fetch0_instr_branch_w = \u_frontend.u_decode.u_dec0.branch_o ;
  assign fetch0_instr_csr_w = \u_frontend.u_decode.u_dec0.csr_o ;
  assign fetch0_instr_div_w = \u_frontend.u_decode.u_dec0.div_o ;
  assign fetch0_instr_exec_w = \u_frontend.u_decode.u_dec0.exec_o ;
  assign fetch0_instr_invalid_w = \u_frontend.u_decode.u_dec0.invalid_w ;
  assign fetch0_instr_lsu_w = \u_frontend.u_decode.u_dec0.lsu_o ;
  assign fetch0_instr_mul_w = \u_frontend.u_decode.u_dec0.mul_o ;
  assign fetch0_instr_rd_valid_w = \u_frontend.u_decode.u_dec0.rd_valid_o ;
  assign fetch0_instr_w = \u_frontend.u_decode.u_fifo.data0_out_o ;
  assign fetch0_pc_w = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h0 };
  assign fetch0_valid_w = \u_frontend.u_decode.u_dec0.valid_i ;
  assign fetch1_accept_w = \u_frontend.u_decode.u_fifo.pop1_i ;
  assign fetch1_fault_fetch_w = \u_frontend.u_decode.u_fifo.info1_out_o [0];
  assign fetch1_fault_page_w = \u_frontend.u_decode.u_fifo.info1_out_o [1];
  assign fetch1_instr_branch_w = \u_frontend.u_decode.u_dec1.branch_o ;
  assign fetch1_instr_csr_w = \u_frontend.u_decode.u_dec1.csr_o ;
  assign fetch1_instr_div_w = \u_frontend.u_decode.u_dec1.div_o ;
  assign fetch1_instr_exec_w = \u_frontend.u_decode.u_dec1.exec_o ;
  assign fetch1_instr_invalid_w = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign fetch1_instr_lsu_w = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign fetch1_instr_mul_w = \u_frontend.u_decode.u_dec1.mul_o ;
  assign fetch1_instr_rd_valid_w = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign fetch1_instr_w = \u_frontend.u_decode.u_fifo.data1_out_o ;
  assign fetch1_pc_w = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign fetch1_valid_w = \u_frontend.u_decode.u_dec1.valid_i ;
  assign ifence_w = \u_csr.ifence_q ;
  assign interrupt_inhibit_w = \u_csr.interrupt_inhibit_i ;
  assign lsu_opcode_opcode_w = \u_issue.lsu_opcode_opcode_o ;
  assign lsu_opcode_ra_operand_w = \u_issue.lsu_opcode_ra_operand_o ;
  assign lsu_opcode_rb_operand_w = \u_issue.lsu_opcode_rb_operand_o ;
  assign lsu_opcode_valid_w = \u_issue.lsu_opcode_valid_o ;
  assign lsu_stall_w = \u_issue.lsu_stall_i ;
  assign mem_d_addr_o = { \u_lsu.mem_addr_q [31:2], 2'h0 };
  assign mem_d_cacheable_o = \u_lsu.mem_cacheable_q ;
  assign mem_d_data_wr_o = \u_lsu.mem_data_wr_q ;
  assign mem_d_flush_o = \u_lsu.mem_flush_q ;
  assign mem_d_invalidate_o = \u_lsu.mem_invalidate_q ;
  assign mem_d_rd_o = \u_lsu.mem_rd_o ;
  assign mem_d_req_tag_o = 11'h000;
  assign mem_d_wr_o = \u_lsu.mem_wr_o ;
  assign mem_d_writeback_o = \u_lsu.mem_writeback_q ;
  assign mem_i_flush_o = \u_frontend.u_fetch.icache_flush_o ;
  assign mem_i_invalidate_o = 1'h0;
  assign mem_i_pc_o = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign mem_i_rd_o = \u_frontend.u_fetch.icache_rd_o ;
  assign mmu_ifetch_accept_w = mem_i_accept_i;
  assign mmu_ifetch_error_w = mem_i_error_i;
  assign mmu_ifetch_flush_w = \u_frontend.u_fetch.icache_flush_o ;
  assign mmu_ifetch_inst_w = mem_i_inst_i;
  assign mmu_ifetch_pc_w = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign mmu_ifetch_rd_w = \u_frontend.u_fetch.icache_rd_o ;
  assign mmu_ifetch_valid_w = mem_i_valid_i;
  assign mmu_lsu_accept_w = mem_d_accept_i;
  assign mmu_lsu_ack_w = mem_d_ack_i;
  assign mmu_lsu_addr_w = { \u_lsu.mem_addr_q [31:2], 2'h0 };
  assign mmu_lsu_cacheable_w = \u_lsu.mem_cacheable_q ;
  assign mmu_lsu_data_rd_w = mem_d_data_rd_i;
  assign mmu_lsu_data_wr_w = \u_lsu.mem_data_wr_q ;
  assign mmu_lsu_error_w = mem_d_error_i;
  assign mmu_lsu_flush_w = \u_lsu.mem_flush_q ;
  assign mmu_lsu_invalidate_w = \u_lsu.mem_invalidate_q ;
  assign mmu_lsu_rd_w = \u_lsu.mem_rd_o ;
  assign mmu_lsu_resp_tag_w = mem_d_resp_tag_i;
  assign mmu_lsu_wr_w = \u_lsu.mem_wr_o ;
  assign mmu_lsu_writeback_w = \u_lsu.mem_writeback_q ;
  assign mmu_mxr_w = \u_csr.u_csrfile.csr_sr_q [19];
  assign mmu_satp_w = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign mmu_sum_w = \u_csr.u_csrfile.csr_sr_q [18];
  assign mul_hold_w = \u_exec0.hold_i ;
  assign mul_opcode_opcode_w = \u_issue.mul_opcode_opcode_o ;
  assign mul_opcode_ra_operand_w = \u_issue.mul_opcode_ra_operand_o ;
  assign mul_opcode_rb_operand_w = \u_issue.mul_opcode_rb_operand_o ;
  assign mul_opcode_valid_w = \u_issue.mul_opcode_valid_o ;
  assign opcode0_opcode_w = \u_csr.opcode_opcode_i ;
  assign opcode0_pc_w = \u_exec0.opcode_pc_i ;
  assign opcode0_ra_idx_w = \u_csr.opcode_opcode_i [19:15];
  assign opcode0_ra_operand_w = \u_csr.opcode_ra_operand_i ;
  assign opcode0_rb_idx_w = \u_csr.opcode_opcode_i [24:20];
  assign opcode0_rb_operand_w = \u_div.opcode_rb_operand_i ;
  assign opcode0_rd_idx_w = \u_csr.opcode_opcode_i [11:7];
  assign opcode1_opcode_w = \u_exec1.opcode_opcode_i ;
  assign opcode1_pc_w = \u_exec1.opcode_pc_i ;
  assign opcode1_ra_idx_w = \u_exec1.opcode_opcode_i [19:15];
  assign opcode1_ra_operand_w = \u_exec1.opcode_ra_operand_i ;
  assign opcode1_rb_idx_w = \u_exec1.opcode_opcode_i [24:20];
  assign opcode1_rb_operand_w = \u_exec1.opcode_rb_operand_i ;
  assign opcode1_rd_idx_w = \u_exec1.opcode_opcode_i [11:7];
  assign take_interrupt_w = \u_csr.take_interrupt_q ;
  assign \u_csr.branch_csr_pc_o = \u_csr.branch_target_q ;
  assign \u_csr.branch_csr_request_o = \u_csr.branch_q ;
  assign \u_csr.clk_i = clk_i;
  assign \u_csr.cpu_id_i = cpu_id_i;
  assign \u_csr.csr_priv_r = \u_csr.opcode_opcode_i [29:28];
  assign \u_csr.csr_result_e1_exception_o = \u_csr.exception_e1_q ;
  assign \u_csr.csr_result_e1_value_o = \u_csr.rd_result_e1_q ;
  assign \u_csr.csr_result_e1_wdata_o = \u_csr.csr_wdata_e1_q ;
  assign \u_csr.csr_result_e1_write_o = \u_csr.rd_valid_e1_q ;
  assign \u_csr.csr_writeback_exception_addr_i = \u_csr.u_csrfile.exception_addr_i ;
  assign \u_csr.csr_writeback_exception_i = \u_csr.u_csrfile.exception_i ;
  assign \u_csr.csr_writeback_exception_pc_i = \u_csr.u_csrfile.exception_pc_i ;
  assign \u_csr.csr_writeback_waddr_i = \u_issue.u_pipe0_ctrl.opcode_wb_q [31:20];
  assign \u_csr.csr_writeback_wdata_i = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  assign \u_csr.csr_writeback_write_i = \u_issue.u_pipe0_ctrl.csr_wr_wb_q ;
  assign \u_csr.current_priv_w = \u_csr.u_csrfile.csr_mpriv_q ;
  assign \u_csr.ifence_o = \u_csr.ifence_q ;
  assign \u_csr.intr_i = intr_i;
  assign \u_csr.mmu_mxr_o = \u_csr.u_csrfile.csr_sr_q [19];
  assign \u_csr.mmu_satp_o = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.mmu_sum_o = \u_csr.u_csrfile.csr_sr_q [18];
  assign \u_csr.opcode_pc_i = \u_exec0.opcode_pc_i ;
  assign \u_csr.opcode_ra_idx_i = \u_csr.opcode_opcode_i [19:15];
  assign \u_csr.opcode_rb_idx_i = \u_csr.opcode_opcode_i [24:20];
  assign \u_csr.opcode_rb_operand_i = \u_div.opcode_rb_operand_i ;
  assign \u_csr.opcode_rd_idx_i = \u_csr.opcode_opcode_i [11:7];
  assign \u_csr.reset_vector_i = reset_vector_i;
  assign \u_csr.rst_i = rst_i;
  assign \u_csr.satp_reg_w = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.status_reg_w = \u_csr.u_csrfile.csr_sr_q ;
  assign \u_csr.take_interrupt_o = \u_csr.take_interrupt_q ;
  assign \u_csr.u_csrfile.branch_r = \u_csr.csr_branch_w ;
  assign \u_csr.u_csrfile.branch_target_r = \u_csr.csr_target_w ;
  assign \u_csr.u_csrfile.clk_i = clk_i;
  assign \u_csr.u_csrfile.cpu_id_i = cpu_id_i;
  assign \u_csr.u_csrfile.csr_branch_o = \u_csr.csr_branch_w ;
  assign \u_csr.u_csrfile.csr_mideleg_q = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.u_csrfile.csr_mip_next_r [31:12] = { \u_csr.u_csrfile.csr_mip_next_q [31:12] };
  assign \u_csr.u_csrfile.csr_mip_next_r [10] = { \u_csr.u_csrfile.csr_mip_next_q [10] };
  assign \u_csr.u_csrfile.csr_mip_next_r [8] = { \u_csr.u_csrfile.csr_mip_next_q [8] };
  assign \u_csr.u_csrfile.csr_mip_next_r [6] = { \u_csr.u_csrfile.csr_mip_next_q [6] };
  assign \u_csr.u_csrfile.csr_mip_next_r [4:0] = { \u_csr.u_csrfile.csr_mip_next_q [4:0] };
  assign \u_csr.u_csrfile.csr_raddr_i = \u_csr.opcode_opcode_i [31:20];
  assign \u_csr.u_csrfile.csr_rdata_o = \u_csr.csr_rdata_w ;
  assign \u_csr.u_csrfile.csr_ren_i = \u_csr.opcode_valid_i ;
  assign \u_csr.u_csrfile.csr_satp_q = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.u_csrfile.csr_sepc_q = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.u_csrfile.csr_stvec_q = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.u_csrfile.csr_target_o = \u_csr.csr_target_w ;
  assign \u_csr.u_csrfile.csr_wdata_i = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  assign \u_csr.u_csrfile.ext_intr_i = intr_i;
  assign \u_csr.u_csrfile.interrupt_o = \u_csr.interrupt_w ;
  assign \u_csr.u_csrfile.irq_masked_r = \u_csr.interrupt_w ;
  assign \u_csr.u_csrfile.priv_o = \u_csr.u_csrfile.csr_mpriv_q ;
  assign \u_csr.u_csrfile.rdata_r = \u_csr.csr_rdata_w ;
  assign \u_csr.u_csrfile.rst_i = rst_i;
  assign \u_csr.u_csrfile.satp_o = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_csr.u_csrfile.status_o = \u_csr.u_csrfile.csr_sr_q ;
  assign \u_div.clk_i = clk_i;
  assign \u_div.opcode_opcode_i = \u_csr.opcode_opcode_i ;
  assign \u_div.opcode_pc_i = \u_exec0.opcode_pc_i ;
  assign \u_div.opcode_ra_idx_i = \u_csr.opcode_opcode_i [19:15];
  assign \u_div.opcode_ra_operand_i = \u_csr.opcode_ra_operand_i ;
  assign \u_div.opcode_rb_idx_i = \u_csr.opcode_opcode_i [24:20];
  assign \u_div.opcode_rd_idx_i = \u_csr.opcode_opcode_i [11:7];
  assign \u_div.rst_i = rst_i;
  assign \u_div.writeback_valid_o = \u_div.valid_q ;
  assign \u_div.writeback_value_o = \u_div.wb_result_q ;
  assign \u_exec0.bimm_r = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [7], \u_csr.opcode_opcode_i [30:25], \u_csr.opcode_opcode_i [11:8], 1'h0 };
  assign \u_exec0.branch_d_pc_o = \u_exec0.branch_target_r ;
  assign \u_exec0.branch_is_call_o = \u_exec0.branch_call_q ;
  assign \u_exec0.branch_is_jmp_o = \u_exec0.branch_jmp_q ;
  assign \u_exec0.branch_is_not_taken_o = \u_exec0.branch_ntaken_q ;
  assign \u_exec0.branch_is_ret_o = \u_exec0.branch_ret_q ;
  assign \u_exec0.branch_is_taken_o = \u_exec0.branch_taken_q ;
  assign \u_exec0.branch_pc_o = \u_exec0.pc_x_q ;
  assign \u_exec0.branch_source_o = \u_exec0.pc_m_q ;
  assign \u_exec0.clk_i = clk_i;
  assign \u_exec0.imm12_r = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31:20] };
  assign \u_exec0.imm20_r = { \u_csr.opcode_opcode_i [31:12], 12'h000 };
  assign \u_exec0.jimm20_r = { \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [31], \u_csr.opcode_opcode_i [19:12], \u_csr.opcode_opcode_i [20], \u_csr.opcode_opcode_i [30:21], 1'h0 };
  assign \u_exec0.opcode_opcode_i = \u_csr.opcode_opcode_i ;
  assign \u_exec0.opcode_ra_idx_i = \u_csr.opcode_opcode_i [19:15];
  assign \u_exec0.opcode_ra_operand_i = \u_csr.opcode_ra_operand_i ;
  assign \u_exec0.opcode_rb_idx_i = \u_csr.opcode_opcode_i [24:20];
  assign \u_exec0.opcode_rb_operand_i = \u_div.opcode_rb_operand_i ;
  assign \u_exec0.opcode_rd_idx_i = \u_csr.opcode_opcode_i [11:7];
  assign \u_exec0.opcode_valid_i = \u_div.opcode_valid_i ;
  assign \u_exec0.rst_i = rst_i;
  assign \u_exec0.shamt_r = \u_csr.opcode_opcode_i [24:20];
  assign \u_exec0.u_alu.alu_a_i = \u_exec0.alu_input_a_r ;
  assign \u_exec0.u_alu.alu_b_i = \u_exec0.alu_input_b_r ;
  assign \u_exec0.u_alu.alu_op_i = \u_exec0.alu_func_r ;
  assign \u_exec0.u_alu.alu_p_o = \u_exec0.alu_p_w ;
  assign \u_exec0.u_alu.result_r = \u_exec0.alu_p_w ;
  assign \u_exec0.writeback_value_o = \u_exec0.result_q ;
  assign \u_exec1.bimm_r = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [7], \u_exec1.opcode_opcode_i [30:25], \u_exec1.opcode_opcode_i [11:8], 1'h0 };
  assign \u_exec1.branch_d_pc_o = \u_exec1.branch_target_r ;
  assign \u_exec1.branch_is_call_o = \u_exec1.branch_call_q ;
  assign \u_exec1.branch_is_jmp_o = \u_exec1.branch_jmp_q ;
  assign \u_exec1.branch_is_not_taken_o = \u_exec1.branch_ntaken_q ;
  assign \u_exec1.branch_is_ret_o = \u_exec1.branch_ret_q ;
  assign \u_exec1.branch_is_taken_o = \u_exec1.branch_taken_q ;
  assign \u_exec1.branch_pc_o = \u_exec1.pc_x_q ;
  assign \u_exec1.branch_source_o = \u_exec1.pc_m_q ;
  assign \u_exec1.clk_i = clk_i;
  assign \u_exec1.hold_i = \u_exec0.hold_i ;
  assign \u_exec1.imm12_r = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31:20] };
  assign \u_exec1.imm20_r = { \u_exec1.opcode_opcode_i [31:12], 12'h000 };
  assign \u_exec1.jimm20_r = { \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [31], \u_exec1.opcode_opcode_i [19:12], \u_exec1.opcode_opcode_i [20], \u_exec1.opcode_opcode_i [30:21], 1'h0 };
  assign \u_exec1.opcode_ra_idx_i = \u_exec1.opcode_opcode_i [19:15];
  assign \u_exec1.opcode_rb_idx_i = \u_exec1.opcode_opcode_i [24:20];
  assign \u_exec1.opcode_rd_idx_i = \u_exec1.opcode_opcode_i [11:7];
  assign \u_exec1.rst_i = rst_i;
  assign \u_exec1.shamt_r = \u_exec1.opcode_opcode_i [24:20];
  assign \u_exec1.u_alu.alu_a_i = \u_exec1.alu_input_a_r ;
  assign \u_exec1.u_alu.alu_b_i = \u_exec1.alu_input_b_r ;
  assign \u_exec1.u_alu.alu_op_i = \u_exec1.alu_func_r ;
  assign \u_exec1.u_alu.alu_p_o = \u_exec1.alu_p_w ;
  assign \u_exec1.u_alu.result_r = \u_exec1.alu_p_w ;
  assign \u_exec1.writeback_value_o = \u_exec1.result_q ;
  assign \u_frontend.branch_info_is_call_i = \u_frontend.u_npc.branch_is_call_i ;
  assign \u_frontend.branch_info_is_jmp_i = \u_frontend.u_npc.branch_is_jmp_i ;
  assign \u_frontend.branch_info_is_not_taken_i = \u_frontend.u_npc.branch_is_not_taken_i ;
  assign \u_frontend.branch_info_is_ret_i = \u_frontend.u_npc.branch_is_ret_i ;
  assign \u_frontend.branch_info_is_taken_i = \u_frontend.u_npc.branch_is_taken_i ;
  assign \u_frontend.branch_info_pc_i = \u_frontend.u_npc.branch_pc_i ;
  assign \u_frontend.branch_info_request_i = \u_frontend.u_npc.branch_request_i ;
  assign \u_frontend.branch_info_source_i = \u_frontend.u_npc.branch_source_i ;
  assign \u_frontend.branch_pc_i = \u_frontend.u_fetch.branch_pc_i ;
  assign \u_frontend.branch_request_i = \u_frontend.u_decode.u_fifo.flush_i ;
  assign \u_frontend.clk_i = clk_i;
  assign \u_frontend.fetch0_accept_i = \u_frontend.u_decode.u_fifo.pop0_i ;
  assign \u_frontend.fetch0_fault_fetch_o = \u_frontend.u_decode.u_fifo.info0_out_o [0];
  assign \u_frontend.fetch0_fault_page_o = \u_frontend.u_decode.u_fifo.info0_out_o [1];
  assign \u_frontend.fetch0_instr_branch_o = \u_frontend.u_decode.u_dec0.branch_o ;
  assign \u_frontend.fetch0_instr_csr_o = \u_frontend.u_decode.u_dec0.csr_o ;
  assign \u_frontend.fetch0_instr_div_o = \u_frontend.u_decode.u_dec0.div_o ;
  assign \u_frontend.fetch0_instr_exec_o = \u_frontend.u_decode.u_dec0.exec_o ;
  assign \u_frontend.fetch0_instr_invalid_o = \u_frontend.u_decode.u_dec0.invalid_w ;
  assign \u_frontend.fetch0_instr_lsu_o = \u_frontend.u_decode.u_dec0.lsu_o ;
  assign \u_frontend.fetch0_instr_mul_o = \u_frontend.u_decode.u_dec0.mul_o ;
  assign \u_frontend.fetch0_instr_o = \u_frontend.u_decode.u_fifo.data0_out_o ;
  assign \u_frontend.fetch0_instr_rd_valid_o = \u_frontend.u_decode.u_dec0.rd_valid_o ;
  assign \u_frontend.fetch0_pc_o = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h0 };
  assign \u_frontend.fetch0_valid_o = \u_frontend.u_decode.u_dec0.valid_i ;
  assign \u_frontend.fetch1_accept_i = \u_frontend.u_decode.u_fifo.pop1_i ;
  assign \u_frontend.fetch1_fault_fetch_o = \u_frontend.u_decode.u_fifo.info1_out_o [0];
  assign \u_frontend.fetch1_fault_page_o = \u_frontend.u_decode.u_fifo.info1_out_o [1];
  assign \u_frontend.fetch1_instr_branch_o = \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_frontend.fetch1_instr_csr_o = \u_frontend.u_decode.u_dec1.csr_o ;
  assign \u_frontend.fetch1_instr_div_o = \u_frontend.u_decode.u_dec1.div_o ;
  assign \u_frontend.fetch1_instr_exec_o = \u_frontend.u_decode.u_dec1.exec_o ;
  assign \u_frontend.fetch1_instr_invalid_o = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_frontend.fetch1_instr_lsu_o = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_frontend.fetch1_instr_mul_o = \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_frontend.fetch1_instr_o = \u_frontend.u_decode.u_fifo.data1_out_o ;
  assign \u_frontend.fetch1_instr_rd_valid_o = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_frontend.fetch1_pc_o = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign \u_frontend.fetch1_valid_o = \u_frontend.u_decode.u_dec1.valid_i ;
  assign \u_frontend.fetch_accept_w = \u_frontend.u_decode.u_fifo.accept_o ;
  assign \u_frontend.fetch_fault_fetch_w = \u_frontend.u_decode.fetch_in_fault_fetch_i ;
  assign \u_frontend.fetch_fault_page_w = \u_frontend.u_decode.fetch_in_fault_page_i ;
  assign \u_frontend.fetch_instr_w = \u_frontend.u_decode.fetch_in_instr_i ;
  assign \u_frontend.fetch_invalidate_i = \u_csr.ifence_q ;
  assign \u_frontend.fetch_pc_accept_w = \u_frontend.u_fetch.pc_accept_o ;
  assign \u_frontend.fetch_pc_f_w = \u_frontend.u_fetch.icache_pc_w ;
  assign \u_frontend.fetch_pc_w = \u_frontend.u_decode.u_fifo.pc_in_i ;
  assign \u_frontend.fetch_pred_branch_w = { \u_frontend.u_fetch.fetch_pred_branch_o [1], \u_frontend.u_decode.u_fifo.pred_in_i [0] };
  assign \u_frontend.fetch_valid_w = \u_frontend.u_decode.u_fifo.push_i ;
  assign \u_frontend.icache_accept_i = mem_i_accept_i;
  assign \u_frontend.icache_error_i = mem_i_error_i;
  assign \u_frontend.icache_flush_o = \u_frontend.u_fetch.icache_flush_o ;
  assign \u_frontend.icache_inst_i = mem_i_inst_i;
  assign \u_frontend.icache_pc_o = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign \u_frontend.icache_rd_o = \u_frontend.u_fetch.icache_rd_o ;
  assign \u_frontend.icache_valid_i = mem_i_valid_i;
  assign \u_frontend.next_pc_f_w = \u_frontend.u_fetch.next_pc_f_i ;
  assign \u_frontend.next_taken_f_w = \u_frontend.u_fetch.next_taken_f_i ;
  assign \u_frontend.rst_i = rst_i;
  assign \u_frontend.u_decode.branch_pc_i = \u_frontend.u_fetch.branch_pc_i ;
  assign \u_frontend.u_decode.branch_request_i = \u_frontend.u_decode.u_fifo.flush_i ;
  assign \u_frontend.u_decode.clk_i = clk_i;
  assign \u_frontend.u_decode.fetch_in_accept_o = \u_frontend.u_decode.u_fifo.accept_o ;
  assign \u_frontend.u_decode.fetch_in_pc_i = \u_frontend.u_decode.u_fifo.pc_in_i ;
  assign \u_frontend.u_decode.fetch_in_pred_branch_i = { \u_frontend.u_fetch.fetch_pred_branch_o [1], \u_frontend.u_decode.u_fifo.pred_in_i [0] };
  assign \u_frontend.u_decode.fetch_in_valid_i = \u_frontend.u_decode.u_fifo.push_i ;
  assign \u_frontend.u_decode.fetch_out0_accept_i = \u_frontend.u_decode.u_fifo.pop0_i ;
  assign \u_frontend.u_decode.fetch_out0_fault_fetch_o = \u_frontend.u_decode.u_fifo.info0_out_o [0];
  assign \u_frontend.u_decode.fetch_out0_fault_page_o = \u_frontend.u_decode.u_fifo.info0_out_o [1];
  assign \u_frontend.u_decode.fetch_out0_instr_branch_o = \u_frontend.u_decode.u_dec0.branch_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_csr_o = \u_frontend.u_decode.u_dec0.csr_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_div_o = \u_frontend.u_decode.u_dec0.div_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_exec_o = \u_frontend.u_decode.u_dec0.exec_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_invalid_o = \u_frontend.u_decode.u_dec0.invalid_w ;
  assign \u_frontend.u_decode.fetch_out0_instr_lsu_o = \u_frontend.u_decode.u_dec0.lsu_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_mul_o = \u_frontend.u_decode.u_dec0.mul_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_o = \u_frontend.u_decode.u_fifo.data0_out_o ;
  assign \u_frontend.u_decode.fetch_out0_instr_rd_valid_o = \u_frontend.u_decode.u_dec0.rd_valid_o ;
  assign \u_frontend.u_decode.fetch_out0_pc_o = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h0 };
  assign \u_frontend.u_decode.fetch_out0_valid_o = \u_frontend.u_decode.u_dec0.valid_i ;
  assign \u_frontend.u_decode.fetch_out1_accept_i = \u_frontend.u_decode.u_fifo.pop1_i ;
  assign \u_frontend.u_decode.fetch_out1_fault_fetch_o = \u_frontend.u_decode.u_fifo.info1_out_o [0];
  assign \u_frontend.u_decode.fetch_out1_fault_page_o = \u_frontend.u_decode.u_fifo.info1_out_o [1];
  assign \u_frontend.u_decode.fetch_out1_instr_branch_o = \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_csr_o = \u_frontend.u_decode.u_dec1.csr_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_div_o = \u_frontend.u_decode.u_dec1.div_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_exec_o = \u_frontend.u_decode.u_dec1.exec_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_invalid_o = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_frontend.u_decode.fetch_out1_instr_lsu_o = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_mul_o = \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_o = \u_frontend.u_decode.u_fifo.data1_out_o ;
  assign \u_frontend.u_decode.fetch_out1_instr_rd_valid_o = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_frontend.u_decode.fetch_out1_pc_o = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign \u_frontend.u_decode.fetch_out1_valid_o = \u_frontend.u_decode.u_dec1.valid_i ;
  assign \u_frontend.u_decode.rst_i = rst_i;
  assign \u_frontend.u_decode.u_dec0.invalid_o = \u_frontend.u_decode.u_dec0.invalid_w ;
  assign \u_frontend.u_decode.u_dec0.opcode_i = \u_frontend.u_decode.u_fifo.data0_out_o ;
  assign \u_frontend.u_decode.u_dec1.invalid_o = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_frontend.u_decode.u_dec1.opcode_i = \u_frontend.u_decode.u_fifo.data1_out_o ;
  assign \u_frontend.u_decode.u_fifo.clk_i = clk_i;
  assign \u_frontend.u_decode.u_fifo.info0_in_i = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign \u_frontend.u_decode.u_fifo.info1_in_i = { \u_frontend.u_decode.fetch_in_fault_page_i , \u_frontend.u_decode.fetch_in_fault_fetch_i };
  assign \u_frontend.u_decode.u_fifo.pc0_out_o [2:0] = 3'h0;
  assign \u_frontend.u_decode.u_fifo.pc1_out_o = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign \u_frontend.u_decode.u_fifo.pred_in_i [1] = \u_frontend.u_fetch.fetch_pred_branch_o [1];
  assign \u_frontend.u_decode.u_fifo.rst_i = rst_i;
  assign \u_frontend.u_decode.u_fifo.valid0_o = \u_frontend.u_decode.u_dec0.valid_i ;
  assign \u_frontend.u_decode.u_fifo.valid1_o = \u_frontend.u_decode.u_dec1.valid_i ;
  assign \u_frontend.u_fetch.branch_request_i = \u_frontend.u_decode.u_fifo.flush_i ;
  assign \u_frontend.u_fetch.clk_i = clk_i;
  assign \u_frontend.u_fetch.fetch_accept_i = \u_frontend.u_decode.u_fifo.accept_o ;
  assign \u_frontend.u_fetch.fetch_fault_fetch_o = \u_frontend.u_decode.fetch_in_fault_fetch_i ;
  assign \u_frontend.u_fetch.fetch_fault_page_o = \u_frontend.u_decode.fetch_in_fault_page_i ;
  assign \u_frontend.u_fetch.fetch_instr_o = \u_frontend.u_decode.fetch_in_instr_i ;
  assign \u_frontend.u_fetch.fetch_invalidate_i = \u_csr.ifence_q ;
  assign \u_frontend.u_fetch.fetch_pc_o = \u_frontend.u_decode.u_fifo.pc_in_i ;
  assign \u_frontend.u_fetch.fetch_pred_branch_o [0] = \u_frontend.u_decode.u_fifo.pred_in_i [0];
  assign \u_frontend.u_fetch.fetch_resp_drop_w = \u_frontend.u_fetch.branch_w ;
  assign \u_frontend.u_fetch.fetch_valid_o = \u_frontend.u_decode.u_fifo.push_i ;
  assign \u_frontend.u_fetch.icache_accept_i = mem_i_accept_i;
  assign \u_frontend.u_fetch.icache_error_i = mem_i_error_i;
  assign \u_frontend.u_fetch.icache_inst_i = mem_i_inst_i;
  assign \u_frontend.u_fetch.icache_pc_o = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign \u_frontend.u_fetch.icache_valid_i = mem_i_valid_i;
  assign \u_frontend.u_fetch.pc_f_o = \u_frontend.u_fetch.icache_pc_w ;
  assign \u_frontend.u_fetch.rst_i = rst_i;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.bht_rd_entry_w = { \u_frontend.u_fetch.icache_pc_w [4:3], \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r };
  assign \u_frontend.u_npc.BRANCH_PREDICTION.bht_wr_entry_w = \u_frontend.u_npc.branch_source_i [4:2];
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_r = \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_call_w ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_r = \u_frontend.u_npc.BRANCH_PREDICTION.btb_is_ret_w ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_w = \u_frontend.u_npc.BRANCH_PREDICTION.btb_upper_r ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_w = \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.btb_wr_alloc_w = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [2:0];
  assign \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.alloc_entry_o = \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.lfsr_q [2:0];
  assign \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.alloc_i = \u_frontend.u_npc.BRANCH_PREDICTION.btb_miss_r ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.clk_i = clk_i;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.hit_i = \u_frontend.u_npc.BRANCH_PREDICTION.btb_valid_r ;
  assign \u_frontend.u_npc.BRANCH_PREDICTION.u_lru.rst_i = rst_i;
  assign \u_frontend.u_npc.clk_i = clk_i;
  assign \u_frontend.u_npc.next_pc_f_o = \u_frontend.u_fetch.next_pc_f_i ;
  assign \u_frontend.u_npc.next_taken_f_o = \u_frontend.u_fetch.next_taken_f_i ;
  assign \u_frontend.u_npc.pc_accept_i = \u_frontend.u_fetch.pc_accept_o ;
  assign \u_frontend.u_npc.pc_f_i = \u_frontend.u_fetch.icache_pc_w ;
  assign \u_frontend.u_npc.rst_i = rst_i;
  assign \u_issue.branch_csr_pc_i = \u_csr.branch_target_q ;
  assign \u_issue.branch_csr_request_i = \u_csr.branch_q ;
  assign \u_issue.branch_d_exec0_pc_i = \u_exec0.branch_target_r ;
  assign \u_issue.branch_d_exec0_request_i = \u_exec0.branch_d_request_o ;
  assign \u_issue.branch_d_exec1_pc_i = \u_exec1.branch_target_r ;
  assign \u_issue.branch_d_exec1_request_i = \u_exec1.branch_d_request_o ;
  assign \u_issue.branch_exec0_is_call_i = \u_exec0.branch_call_q ;
  assign \u_issue.branch_exec0_is_jmp_i = \u_exec0.branch_jmp_q ;
  assign \u_issue.branch_exec0_is_not_taken_i = \u_exec0.branch_ntaken_q ;
  assign \u_issue.branch_exec0_is_ret_i = \u_exec0.branch_ret_q ;
  assign \u_issue.branch_exec0_is_taken_i = \u_exec0.branch_taken_q ;
  assign \u_issue.branch_exec0_pc_i = \u_exec0.pc_x_q ;
  assign \u_issue.branch_exec0_source_i = \u_exec0.pc_m_q ;
  assign \u_issue.branch_exec1_is_call_i = \u_exec1.branch_call_q ;
  assign \u_issue.branch_exec1_is_jmp_i = \u_exec1.branch_jmp_q ;
  assign \u_issue.branch_exec1_is_not_taken_i = \u_exec1.branch_ntaken_q ;
  assign \u_issue.branch_exec1_is_ret_i = \u_exec1.branch_ret_q ;
  assign \u_issue.branch_exec1_is_taken_i = \u_exec1.branch_taken_q ;
  assign \u_issue.branch_exec1_pc_i = \u_exec1.pc_x_q ;
  assign \u_issue.branch_exec1_request_i = \u_exec1.branch_request_o ;
  assign \u_issue.branch_exec1_source_i = \u_exec1.pc_m_q ;
  assign \u_issue.branch_info_is_call_o = \u_frontend.u_npc.branch_is_call_i ;
  assign \u_issue.branch_info_is_jmp_o = \u_frontend.u_npc.branch_is_jmp_i ;
  assign \u_issue.branch_info_is_not_taken_o = \u_frontend.u_npc.branch_is_not_taken_i ;
  assign \u_issue.branch_info_is_ret_o = \u_frontend.u_npc.branch_is_ret_i ;
  assign \u_issue.branch_info_is_taken_o = \u_frontend.u_npc.branch_is_taken_i ;
  assign \u_issue.branch_info_pc_o = \u_frontend.u_npc.branch_pc_i ;
  assign \u_issue.branch_info_request_o = \u_frontend.u_npc.branch_request_i ;
  assign \u_issue.branch_info_source_o = \u_frontend.u_npc.branch_source_i ;
  assign \u_issue.branch_pc_o = \u_frontend.u_fetch.branch_pc_i ;
  assign \u_issue.branch_request_o = \u_frontend.u_decode.u_fifo.flush_i ;
  assign \u_issue.clk_i = clk_i;
  assign \u_issue.csr_opcode_invalid_o = \u_csr.opcode_invalid_i ;
  assign \u_issue.csr_opcode_opcode_o = \u_csr.opcode_opcode_i ;
  assign \u_issue.csr_opcode_pc_o = \u_exec0.opcode_pc_i ;
  assign \u_issue.csr_opcode_ra_idx_o = \u_csr.opcode_opcode_i [19:15];
  assign \u_issue.csr_opcode_ra_operand_o = \u_csr.opcode_ra_operand_i ;
  assign \u_issue.csr_opcode_rb_idx_o = \u_csr.opcode_opcode_i [24:20];
  assign \u_issue.csr_opcode_rb_operand_o = \u_div.opcode_rb_operand_i ;
  assign \u_issue.csr_opcode_rd_idx_o = \u_csr.opcode_opcode_i [11:7];
  assign \u_issue.csr_opcode_valid_o = \u_csr.opcode_valid_i ;
  assign \u_issue.csr_result_e1_exception_i = \u_csr.exception_e1_q ;
  assign \u_issue.csr_result_e1_value_i = \u_csr.rd_result_e1_q ;
  assign \u_issue.csr_result_e1_wdata_i = \u_csr.csr_wdata_e1_q ;
  assign \u_issue.csr_result_e1_write_i = \u_csr.rd_valid_e1_q ;
  assign \u_issue.csr_writeback_exception_addr_o = \u_csr.u_csrfile.exception_addr_i ;
  assign \u_issue.csr_writeback_exception_o = \u_csr.u_csrfile.exception_i ;
  assign \u_issue.csr_writeback_exception_pc_o = \u_csr.u_csrfile.exception_pc_i ;
  assign \u_issue.csr_writeback_waddr_o = \u_issue.u_pipe0_ctrl.opcode_wb_q [31:20];
  assign \u_issue.csr_writeback_wdata_o = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  assign \u_issue.csr_writeback_write_o = \u_issue.u_pipe0_ctrl.csr_wr_wb_q ;
  assign \u_issue.div_opcode_valid_o = \u_div.opcode_valid_i ;
  assign \u_issue.exec0_hold_o = \u_exec0.hold_i ;
  assign \u_issue.exec0_opcode_valid_o = \u_div.opcode_valid_i ;
  assign \u_issue.exec1_hold_o = \u_exec0.hold_i ;
  assign \u_issue.exec1_opcode_valid_o = \u_exec1.opcode_valid_i ;
  assign \u_issue.fetch0_accept_o = \u_frontend.u_decode.u_fifo.pop0_i ;
  assign \u_issue.fetch0_fault_fetch_i = \u_frontend.u_decode.u_fifo.info0_out_o [0];
  assign \u_issue.fetch0_fault_page_i = \u_frontend.u_decode.u_fifo.info0_out_o [1];
  assign \u_issue.fetch0_instr_branch_i = \u_frontend.u_decode.u_dec0.branch_o ;
  assign \u_issue.fetch0_instr_csr_i = \u_frontend.u_decode.u_dec0.csr_o ;
  assign \u_issue.fetch0_instr_div_i = \u_frontend.u_decode.u_dec0.div_o ;
  assign \u_issue.fetch0_instr_exec_i = \u_frontend.u_decode.u_dec0.exec_o ;
  assign \u_issue.fetch0_instr_i = \u_frontend.u_decode.u_fifo.data0_out_o ;
  assign \u_issue.fetch0_instr_invalid_i = \u_frontend.u_decode.u_dec0.invalid_w ;
  assign \u_issue.fetch0_instr_lsu_i = \u_frontend.u_decode.u_dec0.lsu_o ;
  assign \u_issue.fetch0_instr_mul_i = \u_frontend.u_decode.u_dec0.mul_o ;
  assign \u_issue.fetch0_instr_rd_valid_i = \u_frontend.u_decode.u_dec0.rd_valid_o ;
  assign \u_issue.fetch0_pc_i = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h0 };
  assign \u_issue.fetch0_valid_i = \u_frontend.u_decode.u_dec0.valid_i ;
  assign \u_issue.fetch1_accept_o = \u_frontend.u_decode.u_fifo.pop1_i ;
  assign \u_issue.fetch1_fault_fetch_i = \u_frontend.u_decode.u_fifo.info1_out_o [0];
  assign \u_issue.fetch1_fault_page_i = \u_frontend.u_decode.u_fifo.info1_out_o [1];
  assign \u_issue.fetch1_instr_branch_i = \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_issue.fetch1_instr_csr_i = \u_frontend.u_decode.u_dec1.csr_o ;
  assign \u_issue.fetch1_instr_div_i = \u_frontend.u_decode.u_dec1.div_o ;
  assign \u_issue.fetch1_instr_exec_i = \u_frontend.u_decode.u_dec1.exec_o ;
  assign \u_issue.fetch1_instr_i = \u_frontend.u_decode.u_fifo.data1_out_o ;
  assign \u_issue.fetch1_instr_invalid_i = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_issue.fetch1_instr_lsu_i = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_issue.fetch1_instr_mul_i = \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_issue.fetch1_instr_rd_valid_i = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_issue.fetch1_pc_i = { \u_frontend.u_decode.u_fifo.pc0_out_o [31:3], 3'h4 };
  assign \u_issue.fetch1_valid_i = \u_frontend.u_decode.u_dec1.valid_i ;
  assign \u_issue.interrupt_inhibit_o = \u_csr.interrupt_inhibit_i ;
  assign \u_issue.issue_a_ra_idx_w = \u_csr.opcode_opcode_i [19:15];
  assign \u_issue.issue_a_ra_value_r = \u_csr.opcode_ra_operand_i ;
  assign \u_issue.issue_a_rb_idx_w = \u_csr.opcode_opcode_i [24:20];
  assign \u_issue.issue_a_rb_value_r = \u_div.opcode_rb_operand_i ;
  assign \u_issue.issue_a_rd_idx_w = \u_csr.opcode_opcode_i [11:7];
  assign \u_issue.issue_b_branch_w = \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_issue.issue_b_csr_w = \u_frontend.u_decode.u_dec1.csr_o ;
  assign \u_issue.issue_b_div_w = \u_frontend.u_decode.u_dec1.div_o ;
  assign \u_issue.issue_b_exec_w = \u_frontend.u_decode.u_dec1.exec_o ;
  assign \u_issue.issue_b_invalid_w = \u_frontend.u_decode.u_dec1.invalid_w ;
  assign \u_issue.issue_b_lsu_w = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_issue.issue_b_mul_w = \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_issue.issue_b_ra_idx_w = \u_exec1.opcode_opcode_i [19:15];
  assign \u_issue.issue_b_ra_value_r = \u_exec1.opcode_ra_operand_i ;
  assign \u_issue.issue_b_rb_idx_w = \u_exec1.opcode_opcode_i [24:20];
  assign \u_issue.issue_b_rb_value_r = \u_exec1.opcode_rb_operand_i ;
  assign \u_issue.issue_b_rd_idx_w = \u_exec1.opcode_opcode_i [11:7];
  assign \u_issue.issue_b_sb_alloc_w = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_issue.mispredicted_r = \u_frontend.u_npc.branch_request_i ;
  assign \u_issue.mul_hold_o = \u_exec0.hold_i ;
  assign \u_issue.opcode0_opcode_o = \u_csr.opcode_opcode_i ;
  assign \u_issue.opcode0_pc_o = \u_exec0.opcode_pc_i ;
  assign \u_issue.opcode0_ra_idx_o = \u_csr.opcode_opcode_i [19:15];
  assign \u_issue.opcode0_ra_operand_o = \u_csr.opcode_ra_operand_i ;
  assign \u_issue.opcode0_rb_idx_o = \u_csr.opcode_opcode_i [24:20];
  assign \u_issue.opcode0_rb_operand_o = \u_div.opcode_rb_operand_i ;
  assign \u_issue.opcode0_rd_idx_o = \u_csr.opcode_opcode_i [11:7];
  assign \u_issue.opcode1_opcode_o = \u_exec1.opcode_opcode_i ;
  assign \u_issue.opcode1_pc_o = \u_exec1.opcode_pc_i ;
  assign \u_issue.opcode1_ra_idx_o = \u_exec1.opcode_opcode_i [19:15];
  assign \u_issue.opcode1_ra_operand_o = \u_exec1.opcode_ra_operand_i ;
  assign \u_issue.opcode1_rb_idx_o = \u_exec1.opcode_opcode_i [24:20];
  assign \u_issue.opcode1_rb_operand_o = \u_exec1.opcode_rb_operand_i ;
  assign \u_issue.opcode1_rd_idx_o = \u_exec1.opcode_opcode_i [11:7];
  assign \u_issue.opcode_a_accept_r = \u_div.opcode_valid_i ;
  assign \u_issue.opcode_a_issue_r = \u_div.opcode_valid_i ;
  assign \u_issue.opcode_a_pc_r = \u_exec0.opcode_pc_i ;
  assign \u_issue.opcode_a_r = \u_csr.opcode_opcode_i ;
  assign \u_issue.opcode_b_accept_r = \u_exec1.opcode_valid_i ;
  assign \u_issue.opcode_b_issue_r = \u_exec1.opcode_valid_i ;
  assign \u_issue.opcode_b_pc_r = \u_exec1.opcode_pc_i ;
  assign \u_issue.opcode_b_r = \u_exec1.opcode_opcode_i ;
  assign \u_issue.pipe0_branch_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6];
  assign \u_issue.pipe0_exception_wb_w = \u_issue.u_pipe0_ctrl.exception_wb_q ;
  assign \u_issue.pipe0_load_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [1];
  assign \u_issue.pipe0_load_e2_w = \u_issue.u_pipe0_ctrl.ctrl_e2_q [1];
  assign \u_issue.pipe0_mul_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [5];
  assign \u_issue.pipe0_mul_e2_w = \u_issue.u_pipe0_ctrl.ctrl_e2_q [5];
  assign \u_issue.pipe0_opc_wb_w = \u_issue.u_pipe0_ctrl.opcode_wb_q ;
  assign \u_issue.pipe0_opcode_e1_w = \u_issue.u_pipe0_ctrl.opcode_e1_q ;
  assign \u_issue.pipe0_pc_e1_w = \u_issue.u_pipe0_ctrl.pc_e1_q ;
  assign \u_issue.pipe0_pc_wb_w = \u_issue.u_pipe0_ctrl.pc_wb_q ;
  assign \u_issue.pipe0_result_wb_w = \u_issue.u_pipe0_ctrl.result_wb_q ;
  assign \u_issue.pipe0_store_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [2];
  assign \u_issue.pipe0_valid_wb_w = \u_issue.u_pipe0_ctrl.valid_wb_o ;
  assign \u_issue.pipe1_branch_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6];
  assign \u_issue.pipe1_exception_wb_w = \u_issue.u_pipe1_ctrl.exception_wb_q ;
  assign \u_issue.pipe1_load_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [1];
  assign \u_issue.pipe1_load_e2_w = \u_issue.u_pipe1_ctrl.ctrl_e2_q [1];
  assign \u_issue.pipe1_mul_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [5];
  assign \u_issue.pipe1_mul_e2_w = \u_issue.u_pipe1_ctrl.ctrl_e2_q [5];
  assign \u_issue.pipe1_opc_wb_w = \u_issue.u_pipe1_ctrl.opcode_wb_q ;
  assign \u_issue.pipe1_opcode_e1_w = \u_issue.u_pipe1_ctrl.opcode_e1_q ;
  assign \u_issue.pipe1_pc_e1_w = \u_issue.u_pipe1_ctrl.pc_e1_q ;
  assign \u_issue.pipe1_pc_wb_w = \u_issue.u_pipe1_ctrl.pc_wb_q ;
  assign \u_issue.pipe1_result_wb_w = \u_issue.u_pipe1_ctrl.result_wb_q ;
  assign \u_issue.pipe1_store_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [2];
  assign \u_issue.pipe1_valid_wb_w = \u_issue.u_pipe1_ctrl.valid_wb_o ;
  assign \u_issue.rst_i = rst_i;
  assign \u_issue.stall_w = \u_exec0.hold_i ;
  assign \u_issue.take_interrupt_i = \u_csr.take_interrupt_q ;
  assign \u_issue.u_pipe0_ctrl.alu_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [0];
  assign \u_issue.u_pipe0_ctrl.alu_result_e1_i = \u_exec0.result_q ;
  assign \u_issue.u_pipe0_ctrl.branch_e1_o = \u_issue.u_pipe0_ctrl.ctrl_e1_q [6];
  assign \u_issue.u_pipe0_ctrl.clk_i = clk_i;
  assign \u_issue.u_pipe0_ctrl.csr_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [3];
  assign \u_issue.u_pipe0_ctrl.csr_result_exception_e1_i = \u_csr.exception_e1_q ;
  assign \u_issue.u_pipe0_ctrl.csr_result_value_e1_i = \u_csr.rd_result_e1_q ;
  assign \u_issue.u_pipe0_ctrl.csr_result_wdata_e1_i = \u_csr.csr_wdata_e1_q ;
  assign \u_issue.u_pipe0_ctrl.csr_result_write_e1_i = \u_csr.rd_valid_e1_q ;
  assign \u_issue.u_pipe0_ctrl.csr_waddr_wb_o = \u_issue.u_pipe0_ctrl.opcode_wb_q [31:20];
  assign \u_issue.u_pipe0_ctrl.csr_wb_o = \u_issue.pipe0_csr_wb_w ;
  assign \u_issue.u_pipe0_ctrl.csr_wdata_wb_o = \u_issue.u_pipe0_ctrl.csr_wdata_wb_q ;
  assign \u_issue.u_pipe0_ctrl.csr_write_wb_o = \u_issue.u_pipe0_ctrl.csr_wr_wb_q ;
  assign \u_issue.u_pipe0_ctrl.div_complete_i = \u_div.valid_q ;
  assign \u_issue.u_pipe0_ctrl.div_e1_w = \u_issue.u_pipe0_ctrl.ctrl_e1_q [4];
  assign \u_issue.u_pipe0_ctrl.div_result_i = \u_div.wb_result_q ;
  assign \u_issue.u_pipe0_ctrl.exception_wb_o = \u_issue.u_pipe0_ctrl.exception_wb_q ;
  assign \u_issue.u_pipe0_ctrl.issue_accept_i = \u_div.opcode_valid_i ;
  assign \u_issue.u_pipe0_ctrl.issue_branch_i = \u_issue.issue_a_branch_w ;
  assign \u_issue.u_pipe0_ctrl.issue_branch_taken_i = \u_exec0.branch_d_request_o ;
  assign \u_issue.u_pipe0_ctrl.issue_branch_target_i = \u_exec0.branch_target_r ;
  assign \u_issue.u_pipe0_ctrl.issue_csr_i = \u_issue.issue_a_csr_w ;
  assign \u_issue.u_pipe0_ctrl.issue_div_i = \u_issue.issue_a_div_w ;
  assign \u_issue.u_pipe0_ctrl.issue_exception_i = { 1'h0, \u_issue.issue_a_fault_w };
  assign \u_issue.u_pipe0_ctrl.issue_lsu_i = \u_issue.issue_a_lsu_w ;
  assign \u_issue.u_pipe0_ctrl.issue_mul_i = \u_issue.issue_a_mul_w ;
  assign \u_issue.u_pipe0_ctrl.issue_opcode_i = \u_csr.opcode_opcode_i ;
  assign \u_issue.u_pipe0_ctrl.issue_operand_ra_i = \u_csr.opcode_ra_operand_i ;
  assign \u_issue.u_pipe0_ctrl.issue_operand_rb_i = \u_div.opcode_rb_operand_i ;
  assign \u_issue.u_pipe0_ctrl.issue_pc_i = \u_exec0.opcode_pc_i ;
  assign \u_issue.u_pipe0_ctrl.issue_rd_i = \u_csr.opcode_opcode_i [11:7];
  assign \u_issue.u_pipe0_ctrl.issue_rd_valid_i = \u_issue.issue_a_sb_alloc_w ;
  assign \u_issue.u_pipe0_ctrl.issue_stall_i = \u_exec0.hold_i ;
  assign \u_issue.u_pipe0_ctrl.issue_valid_i = \u_div.opcode_valid_i ;
  assign \u_issue.u_pipe0_ctrl.load_e1_o = \u_issue.u_pipe0_ctrl.ctrl_e1_q [1];
  assign \u_issue.u_pipe0_ctrl.load_e2_o = \u_issue.u_pipe0_ctrl.ctrl_e2_q [1];
  assign \u_issue.u_pipe0_ctrl.mem_exception_e2_i [5] = 1'h0;
  assign \u_issue.u_pipe0_ctrl.mul_e1_o = \u_issue.u_pipe0_ctrl.ctrl_e1_q [5];
  assign \u_issue.u_pipe0_ctrl.mul_e2_o = \u_issue.u_pipe0_ctrl.ctrl_e2_q [5];
  assign \u_issue.u_pipe0_ctrl.mul_result_e2_i = \u_mul.result_e2_q ;
  assign \u_issue.u_pipe0_ctrl.opcode_e1_o = \u_issue.u_pipe0_ctrl.opcode_e1_q ;
  assign \u_issue.u_pipe0_ctrl.opcode_wb_o = \u_issue.u_pipe0_ctrl.opcode_wb_q ;
  assign \u_issue.u_pipe0_ctrl.pc_e1_o = \u_issue.u_pipe0_ctrl.pc_e1_q ;
  assign \u_issue.u_pipe0_ctrl.pc_wb_o = \u_issue.u_pipe0_ctrl.pc_wb_q ;
  assign \u_issue.u_pipe0_ctrl.rd_e1_o = \u_issue.pipe0_rd_e1_w ;
  assign \u_issue.u_pipe0_ctrl.rd_e2_o = \u_issue.pipe0_rd_e2_w ;
  assign \u_issue.u_pipe0_ctrl.rd_wb_o = \u_issue.pipe0_rd_wb_w ;
  assign \u_issue.u_pipe0_ctrl.result_e2_o = \u_issue.pipe0_result_e2_w ;
  assign \u_issue.u_pipe0_ctrl.result_e2_r = \u_issue.pipe0_result_e2_w ;
  assign \u_issue.u_pipe0_ctrl.result_wb_o = \u_issue.u_pipe0_ctrl.result_wb_q ;
  assign \u_issue.u_pipe0_ctrl.rst_i = rst_i;
  assign \u_issue.u_pipe0_ctrl.squash_e1_e2_i = \u_issue.pipe1_squash_e1_e2_w ;
  assign \u_issue.u_pipe0_ctrl.squash_e1_e2_o = \u_issue.pipe0_squash_e1_e2_w ;
  assign \u_issue.u_pipe0_ctrl.stall_o = \u_issue.pipe0_stall_raw_w ;
  assign \u_issue.u_pipe0_ctrl.store_e1_o = \u_issue.u_pipe0_ctrl.ctrl_e1_q [2];
  assign \u_issue.u_pipe0_ctrl.take_interrupt_i = \u_csr.take_interrupt_q ;
  assign \u_issue.u_pipe1_ctrl.alu_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [0];
  assign \u_issue.u_pipe1_ctrl.alu_result_e1_i = \u_exec1.result_q ;
  assign \u_issue.u_pipe1_ctrl.branch_e1_o = \u_issue.u_pipe1_ctrl.ctrl_e1_q [6];
  assign \u_issue.u_pipe1_ctrl.clk_i = clk_i;
  assign \u_issue.u_pipe1_ctrl.csr_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [3];
  assign \u_issue.u_pipe1_ctrl.csr_result_exception_e1_i = \u_csr.exception_e1_q ;
  assign \u_issue.u_pipe1_ctrl.csr_result_value_e1_i = \u_csr.rd_result_e1_q ;
  assign \u_issue.u_pipe1_ctrl.csr_result_wdata_e1_i = \u_csr.csr_wdata_e1_q ;
  assign \u_issue.u_pipe1_ctrl.csr_result_write_e1_i = \u_csr.rd_valid_e1_q ;
  assign \u_issue.u_pipe1_ctrl.csr_waddr_wb_o = \u_issue.u_pipe1_ctrl.opcode_wb_q [31:20];
  assign \u_issue.u_pipe1_ctrl.div_complete_i = \u_div.valid_q ;
  assign \u_issue.u_pipe1_ctrl.div_e1_w = \u_issue.u_pipe1_ctrl.ctrl_e1_q [4];
  assign \u_issue.u_pipe1_ctrl.div_result_i = \u_div.wb_result_q ;
  assign \u_issue.u_pipe1_ctrl.exception_wb_o = \u_issue.u_pipe1_ctrl.exception_wb_q ;
  assign \u_issue.u_pipe1_ctrl.issue_accept_i = \u_exec1.opcode_valid_i ;
  assign \u_issue.u_pipe1_ctrl.issue_branch_i = \u_frontend.u_decode.u_dec1.branch_o ;
  assign \u_issue.u_pipe1_ctrl.issue_branch_taken_i = \u_exec1.branch_d_request_o ;
  assign \u_issue.u_pipe1_ctrl.issue_branch_target_i = \u_exec1.branch_target_r ;
  assign \u_issue.u_pipe1_ctrl.issue_exception_i = { 1'h0, \u_issue.issue_b_fault_w };
  assign \u_issue.u_pipe1_ctrl.issue_lsu_i = \u_frontend.u_decode.u_dec1.lsu_o ;
  assign \u_issue.u_pipe1_ctrl.issue_mul_i = \u_frontend.u_decode.u_dec1.mul_o ;
  assign \u_issue.u_pipe1_ctrl.issue_opcode_i = \u_exec1.opcode_opcode_i ;
  assign \u_issue.u_pipe1_ctrl.issue_operand_ra_i = \u_exec1.opcode_ra_operand_i ;
  assign \u_issue.u_pipe1_ctrl.issue_operand_rb_i = \u_exec1.opcode_rb_operand_i ;
  assign \u_issue.u_pipe1_ctrl.issue_pc_i = \u_exec1.opcode_pc_i ;
  assign \u_issue.u_pipe1_ctrl.issue_rd_i = \u_exec1.opcode_opcode_i [11:7];
  assign \u_issue.u_pipe1_ctrl.issue_rd_valid_i = \u_frontend.u_decode.u_dec1.rd_valid_o ;
  assign \u_issue.u_pipe1_ctrl.issue_stall_i = \u_exec0.hold_i ;
  assign \u_issue.u_pipe1_ctrl.issue_valid_i = \u_exec1.opcode_valid_i ;
  assign \u_issue.u_pipe1_ctrl.load_e1_o = \u_issue.u_pipe1_ctrl.ctrl_e1_q [1];
  assign \u_issue.u_pipe1_ctrl.load_e2_o = \u_issue.u_pipe1_ctrl.ctrl_e2_q [1];
  assign \u_issue.u_pipe1_ctrl.mem_complete_i = \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign \u_issue.u_pipe1_ctrl.mem_exception_e2_i = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign \u_issue.u_pipe1_ctrl.mem_result_e2_i = \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  assign \u_issue.u_pipe1_ctrl.mul_e1_o = \u_issue.u_pipe1_ctrl.ctrl_e1_q [5];
  assign \u_issue.u_pipe1_ctrl.mul_e2_o = \u_issue.u_pipe1_ctrl.ctrl_e2_q [5];
  assign \u_issue.u_pipe1_ctrl.mul_result_e2_i = \u_mul.result_e2_q ;
  assign \u_issue.u_pipe1_ctrl.opcode_e1_o = \u_issue.u_pipe1_ctrl.opcode_e1_q ;
  assign \u_issue.u_pipe1_ctrl.opcode_wb_o = \u_issue.u_pipe1_ctrl.opcode_wb_q ;
  assign \u_issue.u_pipe1_ctrl.pc_e1_o = \u_issue.u_pipe1_ctrl.pc_e1_q ;
  assign \u_issue.u_pipe1_ctrl.pc_wb_o = \u_issue.u_pipe1_ctrl.pc_wb_q ;
  assign \u_issue.u_pipe1_ctrl.rd_e1_o = \u_issue.pipe1_rd_e1_w ;
  assign \u_issue.u_pipe1_ctrl.rd_e2_o = \u_issue.pipe1_rd_e2_w ;
  assign \u_issue.u_pipe1_ctrl.rd_wb_o = \u_issue.pipe1_rd_wb_w ;
  assign \u_issue.u_pipe1_ctrl.result_e2_o = \u_issue.pipe1_result_e2_w ;
  assign \u_issue.u_pipe1_ctrl.result_e2_r = \u_issue.pipe1_result_e2_w ;
  assign \u_issue.u_pipe1_ctrl.result_wb_o = \u_issue.u_pipe1_ctrl.result_wb_q ;
  assign \u_issue.u_pipe1_ctrl.rst_i = rst_i;
  assign \u_issue.u_pipe1_ctrl.squash_e1_e2_i = \u_issue.pipe0_squash_e1_e2_w ;
  assign \u_issue.u_pipe1_ctrl.squash_e1_e2_o = \u_issue.pipe1_squash_e1_e2_w ;
  assign \u_issue.u_pipe1_ctrl.squash_wb_i = \u_issue.pipe0_squash_e1_e2_w ;
  assign \u_issue.u_pipe1_ctrl.stall_o = \u_issue.pipe1_stall_raw_w ;
  assign \u_issue.u_pipe1_ctrl.store_e1_o = \u_issue.u_pipe1_ctrl.ctrl_e1_q [2];
  assign \u_issue.u_pipe1_ctrl.take_interrupt_i = \u_csr.take_interrupt_q ;
  assign \u_issue.u_regfile.REGFILE.ra0_value_r = \u_issue.issue_a_ra_value_w ;
  assign \u_issue.u_regfile.REGFILE.ra1_value_r = \u_issue.issue_b_ra_value_w ;
  assign \u_issue.u_regfile.REGFILE.rb0_value_r = \u_issue.issue_a_rb_value_w ;
  assign \u_issue.u_regfile.REGFILE.rb1_value_r = \u_issue.issue_b_rb_value_w ;
  assign \u_issue.u_regfile.REGFILE.x10_a0_w = \u_issue.u_regfile.REGFILE.reg_r10_q ;
  assign \u_issue.u_regfile.REGFILE.x11_a1_w = \u_issue.u_regfile.REGFILE.reg_r11_q ;
  assign \u_issue.u_regfile.REGFILE.x12_a2_w = \u_issue.u_regfile.REGFILE.reg_r12_q ;
  assign \u_issue.u_regfile.REGFILE.x13_a3_w = \u_issue.u_regfile.REGFILE.reg_r13_q ;
  assign \u_issue.u_regfile.REGFILE.x14_a4_w = \u_issue.u_regfile.REGFILE.reg_r14_q ;
  assign \u_issue.u_regfile.REGFILE.x15_a5_w = \u_issue.u_regfile.REGFILE.reg_r15_q ;
  assign \u_issue.u_regfile.REGFILE.x16_a6_w = \u_issue.u_regfile.REGFILE.reg_r16_q ;
  assign \u_issue.u_regfile.REGFILE.x17_a7_w = \u_issue.u_regfile.REGFILE.reg_r17_q ;
  assign \u_issue.u_regfile.REGFILE.x18_s2_w = \u_issue.u_regfile.REGFILE.reg_r18_q ;
  assign \u_issue.u_regfile.REGFILE.x19_s3_w = \u_issue.u_regfile.REGFILE.reg_r19_q ;
  assign \u_issue.u_regfile.REGFILE.x1_ra_w = \u_issue.u_regfile.REGFILE.reg_r1_q ;
  assign \u_issue.u_regfile.REGFILE.x20_s4_w = \u_issue.u_regfile.REGFILE.reg_r20_q ;
  assign \u_issue.u_regfile.REGFILE.x21_s5_w = \u_issue.u_regfile.REGFILE.reg_r21_q ;
  assign \u_issue.u_regfile.REGFILE.x22_s6_w = \u_issue.u_regfile.REGFILE.reg_r22_q ;
  assign \u_issue.u_regfile.REGFILE.x23_s7_w = \u_issue.u_regfile.REGFILE.reg_r23_q ;
  assign \u_issue.u_regfile.REGFILE.x24_s8_w = \u_issue.u_regfile.REGFILE.reg_r24_q ;
  assign \u_issue.u_regfile.REGFILE.x25_s9_w = \u_issue.u_regfile.REGFILE.reg_r25_q ;
  assign \u_issue.u_regfile.REGFILE.x26_s10_w = \u_issue.u_regfile.REGFILE.reg_r26_q ;
  assign \u_issue.u_regfile.REGFILE.x27_s11_w = \u_issue.u_regfile.REGFILE.reg_r27_q ;
  assign \u_issue.u_regfile.REGFILE.x28_t3_w = \u_issue.u_regfile.REGFILE.reg_r28_q ;
  assign \u_issue.u_regfile.REGFILE.x29_t4_w = \u_issue.u_regfile.REGFILE.reg_r29_q ;
  assign \u_issue.u_regfile.REGFILE.x2_sp_w = \u_issue.u_regfile.REGFILE.reg_r2_q ;
  assign \u_issue.u_regfile.REGFILE.x30_t5_w = \u_issue.u_regfile.REGFILE.reg_r30_q ;
  assign \u_issue.u_regfile.REGFILE.x31_t6_w = \u_issue.u_regfile.REGFILE.reg_r31_q ;
  assign \u_issue.u_regfile.REGFILE.x3_gp_w = \u_issue.u_regfile.REGFILE.reg_r3_q ;
  assign \u_issue.u_regfile.REGFILE.x4_tp_w = \u_issue.u_regfile.REGFILE.reg_r4_q ;
  assign \u_issue.u_regfile.REGFILE.x5_t0_w = \u_issue.u_regfile.REGFILE.reg_r5_q ;
  assign \u_issue.u_regfile.REGFILE.x6_t1_w = \u_issue.u_regfile.REGFILE.reg_r6_q ;
  assign \u_issue.u_regfile.REGFILE.x7_t2_w = \u_issue.u_regfile.REGFILE.reg_r7_q ;
  assign \u_issue.u_regfile.REGFILE.x8_s0_w = \u_issue.u_regfile.REGFILE.reg_r8_q ;
  assign \u_issue.u_regfile.REGFILE.x9_s1_w = \u_issue.u_regfile.REGFILE.reg_r9_q ;
  assign \u_issue.u_regfile.clk_i = clk_i;
  assign \u_issue.u_regfile.ra0_i = \u_csr.opcode_opcode_i [19:15];
  assign \u_issue.u_regfile.ra0_value_o = \u_issue.issue_a_ra_value_w ;
  assign \u_issue.u_regfile.ra1_i = \u_exec1.opcode_opcode_i [19:15];
  assign \u_issue.u_regfile.ra1_value_o = \u_issue.issue_b_ra_value_w ;
  assign \u_issue.u_regfile.rb0_i = \u_csr.opcode_opcode_i [24:20];
  assign \u_issue.u_regfile.rb0_value_o = \u_issue.issue_a_rb_value_w ;
  assign \u_issue.u_regfile.rb1_i = \u_exec1.opcode_opcode_i [24:20];
  assign \u_issue.u_regfile.rb1_value_o = \u_issue.issue_b_rb_value_w ;
  assign \u_issue.u_regfile.rd0_i = \u_issue.pipe0_rd_wb_w ;
  assign \u_issue.u_regfile.rd0_value_i = \u_issue.u_pipe0_ctrl.result_wb_q ;
  assign \u_issue.u_regfile.rd1_i = \u_issue.pipe1_rd_wb_w ;
  assign \u_issue.u_regfile.rd1_value_i = \u_issue.u_pipe1_ctrl.result_wb_q ;
  assign \u_issue.u_regfile.rst_i = rst_i;
  assign \u_issue.writeback_div_valid_i = \u_div.valid_q ;
  assign \u_issue.writeback_div_value_i = \u_div.wb_result_q ;
  assign \u_issue.writeback_exec0_value_i = \u_exec0.result_q ;
  assign \u_issue.writeback_exec1_value_i = \u_exec1.result_q ;
  assign \u_issue.writeback_mem_exception_i = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign \u_issue.writeback_mem_valid_i = \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign \u_issue.writeback_mem_value_i = \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  assign \u_issue.writeback_mul_value_i = \u_mul.result_e2_q ;
  assign \u_lsu.addr_lsb_r = \u_lsu.u_lsu_request.data_out_o [5:4];
  assign \u_lsu.clk_i = clk_i;
  assign \u_lsu.load_byte_r = \u_lsu.u_lsu_request.data_out_o [1];
  assign \u_lsu.load_half_r = \u_lsu.u_lsu_request.data_out_o [2];
  assign \u_lsu.load_signed_r = \u_lsu.u_lsu_request.data_out_o [3];
  assign \u_lsu.mem_accept_i = mem_d_accept_i;
  assign \u_lsu.mem_ack_i = mem_d_ack_i;
  assign \u_lsu.mem_addr_o = { \u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u_lsu.mem_cacheable_o = \u_lsu.mem_cacheable_q ;
  assign \u_lsu.mem_data_rd_i = mem_d_data_rd_i;
  assign \u_lsu.mem_data_wr_o = \u_lsu.mem_data_wr_q ;
  assign \u_lsu.mem_error_i = mem_d_error_i;
  assign \u_lsu.mem_flush_o = \u_lsu.mem_flush_q ;
  assign \u_lsu.mem_invalidate_o = \u_lsu.mem_invalidate_q ;
  assign \u_lsu.mem_resp_tag_i = mem_d_resp_tag_i;
  assign \u_lsu.mem_writeback_o = \u_lsu.mem_writeback_q ;
  assign \u_lsu.opcode_opcode_i = \u_issue.lsu_opcode_opcode_o ;
  assign \u_lsu.opcode_ra_operand_i = \u_issue.lsu_opcode_ra_operand_o ;
  assign \u_lsu.opcode_rb_operand_i = \u_issue.lsu_opcode_rb_operand_o ;
  assign \u_lsu.opcode_valid_i = \u_issue.lsu_opcode_valid_o ;
  assign \u_lsu.resp_addr_w = \u_lsu.u_lsu_request.data_out_o [35:4];
  assign \u_lsu.resp_byte_w = \u_lsu.u_lsu_request.data_out_o [1];
  assign \u_lsu.resp_half_w = \u_lsu.u_lsu_request.data_out_o [2];
  assign \u_lsu.resp_load_w = \u_lsu.u_lsu_request.data_out_o [0];
  assign \u_lsu.resp_signed_w = \u_lsu.u_lsu_request.data_out_o [3];
  assign \u_lsu.rst_i = rst_i;
  assign \u_lsu.stall_o = \u_issue.lsu_stall_i ;
  assign \u_lsu.u_lsu_request.clk_i = clk_i;
  assign \u_lsu.u_lsu_request.data_in_i = { \u_lsu.mem_addr_q , \u_lsu.mem_ls_q , \u_lsu.mem_xh_q , \u_lsu.mem_xb_q , \u_lsu.mem_load_q };
  assign \u_lsu.u_lsu_request.rst_i = rst_i;
  assign \u_lsu.wb_result_r = \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  assign \u_lsu.writeback_exception_o = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign \u_lsu.writeback_valid_o = \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign \u_lsu.writeback_value_o = \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  assign \u_mmu.clk_i = clk_i;
  assign \u_mmu.fetch_in_accept_o = mem_i_accept_i;
  assign \u_mmu.fetch_in_error_o = mem_i_error_i;
  assign \u_mmu.fetch_in_flush_i = \u_frontend.u_fetch.icache_flush_o ;
  assign \u_mmu.fetch_in_inst_o = mem_i_inst_i;
  assign \u_mmu.fetch_in_pc_i = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign \u_mmu.fetch_in_rd_i = \u_frontend.u_fetch.icache_rd_o ;
  assign \u_mmu.fetch_in_valid_o = mem_i_valid_i;
  assign \u_mmu.fetch_out_accept_i = mem_i_accept_i;
  assign \u_mmu.fetch_out_error_i = mem_i_error_i;
  assign \u_mmu.fetch_out_flush_o = \u_frontend.u_fetch.icache_flush_o ;
  assign \u_mmu.fetch_out_inst_i = mem_i_inst_i;
  assign \u_mmu.fetch_out_pc_o = { \u_frontend.u_fetch.icache_pc_w [31:3], 3'h0 };
  assign \u_mmu.fetch_out_rd_o = \u_frontend.u_fetch.icache_rd_o ;
  assign \u_mmu.fetch_out_valid_i = mem_i_valid_i;
  assign \u_mmu.lsu_in_accept_o = mem_d_accept_i;
  assign \u_mmu.lsu_in_ack_o = mem_d_ack_i;
  assign \u_mmu.lsu_in_addr_i = { \u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u_mmu.lsu_in_cacheable_i = \u_lsu.mem_cacheable_q ;
  assign \u_mmu.lsu_in_data_rd_o = mem_d_data_rd_i;
  assign \u_mmu.lsu_in_data_wr_i = \u_lsu.mem_data_wr_q ;
  assign \u_mmu.lsu_in_error_o = mem_d_error_i;
  assign \u_mmu.lsu_in_flush_i = \u_lsu.mem_flush_q ;
  assign \u_mmu.lsu_in_invalidate_i = \u_lsu.mem_invalidate_q ;
  assign \u_mmu.lsu_in_rd_i = \u_lsu.mem_rd_o ;
  assign \u_mmu.lsu_in_resp_tag_o = mem_d_resp_tag_i;
  assign \u_mmu.lsu_in_wr_i = \u_lsu.mem_wr_o ;
  assign \u_mmu.lsu_in_writeback_i = \u_lsu.mem_writeback_q ;
  assign \u_mmu.lsu_out_accept_i = mem_d_accept_i;
  assign \u_mmu.lsu_out_ack_i = mem_d_ack_i;
  assign \u_mmu.lsu_out_addr_o = { \u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u_mmu.lsu_out_cacheable_o = \u_lsu.mem_cacheable_q ;
  assign \u_mmu.lsu_out_data_rd_i = mem_d_data_rd_i;
  assign \u_mmu.lsu_out_data_wr_o = \u_lsu.mem_data_wr_q ;
  assign \u_mmu.lsu_out_error_i = mem_d_error_i;
  assign \u_mmu.lsu_out_flush_o = \u_lsu.mem_flush_q ;
  assign \u_mmu.lsu_out_invalidate_o = \u_lsu.mem_invalidate_q ;
  assign \u_mmu.lsu_out_rd_o = \u_lsu.mem_rd_o ;
  assign \u_mmu.lsu_out_resp_tag_i = mem_d_resp_tag_i;
  assign \u_mmu.lsu_out_wr_o = \u_lsu.mem_wr_o ;
  assign \u_mmu.lsu_out_writeback_o = \u_lsu.mem_writeback_q ;
  assign \u_mmu.mxr_i = \u_csr.u_csrfile.csr_sr_q [19];
  assign \u_mmu.rst_i = rst_i;
  assign \u_mmu.satp_i = \u_csr.u_csrfile.csr_mtimecmp_q ;
  assign \u_mmu.sum_i = \u_csr.u_csrfile.csr_sr_q [18];
  assign \u_mul.clk_i = clk_i;
  assign \u_mul.hold_i = \u_exec0.hold_i ;
  assign \u_mul.opcode_opcode_i = \u_issue.mul_opcode_opcode_o ;
  assign \u_mul.opcode_ra_operand_i = \u_issue.mul_opcode_ra_operand_o ;
  assign \u_mul.opcode_rb_operand_i = \u_issue.mul_opcode_rb_operand_o ;
  assign \u_mul.opcode_valid_i = \u_issue.mul_opcode_valid_o ;
  assign \u_mul.rst_i = rst_i;
  assign \u_mul.writeback_value_o = \u_mul.result_e2_q ;
  assign writeback_div_valid_w = \u_div.valid_q ;
  assign writeback_div_value_w = \u_div.wb_result_q ;
  assign writeback_exec0_value_w = \u_exec0.result_q ;
  assign writeback_exec1_value_w = \u_exec1.result_q ;
  assign writeback_mem_exception_w = { 1'h0, \u_issue.u_pipe0_ctrl.mem_exception_e2_i [4:0] };
  assign writeback_mem_valid_w = \u_issue.u_pipe0_ctrl.mem_complete_i ;
  assign writeback_mem_value_w = \u_issue.u_pipe0_ctrl.mem_result_e2_i ;
  assign writeback_mul_value_w = \u_mul.result_e2_q ;
endmodule
