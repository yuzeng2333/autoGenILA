module CDMA_leading_sign_17_0(mantissa, rtn);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:311" *)
  wire _000_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *)
  wire _001_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:319" *)
  wire _002_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *)
  wire _003_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *)
  wire _004_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *)
  wire _005_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _006_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _007_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _008_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _009_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _010_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _011_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *)
  wire _012_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:303" *)
  wire _013_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:310" *)
  wire _014_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:299" *)
  wire _015_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:300" *)
  wire _016_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:301" *)
  wire _017_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:305" *)
  wire _018_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:306" *)
  wire _019_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:307" *)
  wire _020_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *)
  wire _021_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _022_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _023_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _024_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:313" *)
  wire _025_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *)
  wire _026_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *)
  wire _027_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *)
  wire _028_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *)
  wire _029_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *)
  wire _030_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *)
  wire _031_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *)
  wire _032_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _033_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _034_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _035_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _036_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _037_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _038_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _039_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _040_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _041_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *)
  wire _042_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *)
  wire _043_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *)
  wire _044_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:316" *)
  wire _045_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:319" *)
  wire _046_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *)
  wire _047_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *)
  wire _048_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *)
  wire _049_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _050_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *)
  wire _051_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *)
  wire _052_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *)
  wire _053_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:296" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:295" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:297" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:294" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:287" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:283" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:288" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:284" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:289" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:285" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:286" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:282" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:290" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:291" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:292" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:293" *)
  wire c_h_1_7;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:279" *)
  input [16:0] mantissa;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:280" *)
  output [4:0] rtn;
  assign c_h_1_2 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:302" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3 = _013_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:304" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:308" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:309" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _014_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:311" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:311" *) c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:312" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl = c_h_1_6 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:313" *) _025_;
  assign _001_ = c_h_1_2 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *) _044_;
  assign _002_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:319" *) _046_;
  assign _003_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *) _047_;
  assign _004_ = _028_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) c_h_1_6;
  assign _005_ = _002_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) _029_;
  assign _006_ = _050_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) c_h_1_2;
  assign _007_ = _032_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _034_;
  assign _008_ = _052_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) c_h_1_5;
  assign _009_ = _036_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _038_;
  assign _010_ = _039_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) c_h_1_6;
  assign _011_ = _007_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _040_;
  assign _012_ = _043_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *) c_h_1_7;
  assign _013_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:303" *) mantissa[10:9];
  assign _014_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:310" *) mantissa[2:1];
  assign _015_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:299" *) mantissa[14:13];
  assign _016_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:300" *) mantissa[16:15];
  assign _017_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:301" *) mantissa[12:11];
  assign _018_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:305" *) mantissa[6:5];
  assign _019_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:306" *) mantissa[8:7];
  assign _020_ = | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:307" *) mantissa[4:3];
  assign _021_ = mantissa[15:14] != (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *) 1'b1;
  assign _022_ = mantissa[11:10] != (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) 1'b1;
  assign _023_ = mantissa[7:6] != (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) 1'b1;
  assign _024_ = mantissa[3:2] != (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) 1'b1;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:299" *) _015_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:300" *) _016_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:301" *) _017_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:305" *) _018_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:306" *) _019_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:307" *) _020_;
  assign _025_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:313" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  assign _026_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  assign _027_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *) _001_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:316" *) _045_;
  assign _028_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *) _003_;
  assign _029_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) _004_;
  assign _030_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) _005_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) _048_;
  assign _031_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *) _021_;
  assign _032_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *) _049_;
  assign _033_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _022_;
  assign _034_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _006_;
  assign _035_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _023_;
  assign _036_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _051_;
  assign _037_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _024_;
  assign _038_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _008_;
  assign _039_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _009_;
  assign _040_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _010_;
  assign _041_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _011_;
  assign _042_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *) _053_;
  assign _043_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *) mantissa[0];
  assign _044_ = c_h_1_5 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:315" *) _026_;
  assign _045_ = _027_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:316" *) c_h_1_7;
  assign _046_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:319" *) _015_;
  assign _047_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:320" *) _018_;
  assign _048_ = _030_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:321" *) c_h_1_7;
  assign _049_ = mantissa[16] | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:323" *) _031_;
  assign _050_ = mantissa[12] | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _033_;
  assign _051_ = mantissa[8] | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:324" *) _035_;
  assign _052_ = mantissa[4] | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:325" *) _037_;
  assign _053_ = _041_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *) c_h_1_7;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl = _042_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:326" *) _012_;
  assign rtn = { c_h_1_7, IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl };
endmodule
