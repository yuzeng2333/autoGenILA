module NV_NVDLA_MCIF_READ_cq(nvdla_core_clk, nvdla_core_rstn, cq_wr_prdy, cq_wr_pvld, cq_wr_thread_id, cq_wr_pd, cq_rd0_prdy, cq_rd0_pvld, cq_rd0_pd, cq_rd1_prdy, cq_rd1_pvld, cq_rd1_pd, cq_rd2_prdy, cq_rd2_pvld, cq_rd2_pd, cq_rd3_prdy, cq_rd3_pvld, cq_rd3_pd, cq_rd4_prdy, cq_rd4_pvld, cq_rd4_pd, cq_rd5_prdy, cq_rd5_pvld, cq_rd5_pd, cq_rd6_prdy, cq_rd6_pvld, cq_rd6_pd, cq_rd7_prdy, cq_rd7_pvld, cq_rd7_pd, cq_rd8_prdy, cq_rd8_pvld, cq_rd8_pd, cq_rd9_prdy, cq_rd9_pvld, cq_rd9_pd, pwrbus_ram_pd);
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2628" *)
  wire [8:0] _0000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2628" *)
  wire _0001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2724" *)
  wire [8:0] _0002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2724" *)
  wire _0003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2820" *)
  wire [8:0] _0004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2820" *)
  wire _0005_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2916" *)
  wire [8:0] _0006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2916" *)
  wire _0007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3012" *)
  wire [8:0] _0008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3012" *)
  wire _0009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3108" *)
  wire [8:0] _0010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3108" *)
  wire _0011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3204" *)
  wire [8:0] _0012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3204" *)
  wire _0013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3300" *)
  wire [8:0] _0014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3300" *)
  wire _0015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3396" *)
  wire [8:0] _0016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3396" *)
  wire _0017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3492" *)
  wire [8:0] _0018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3492" *)
  wire _0019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2143" *)
  wire [8:0] _0029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2007" *)
  wire [9:0] _0030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3615" *)
  wire [3:0] _0031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:156" *)
  wire [8:0] _0032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:207" *)
  wire [254:0] _0033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2537" *)
  wire [7:0] _0044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2007" *)
  wire _0045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2568" *)
  wire [6:0] _0046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2603" *)
  wire _0047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2568" *)
  wire [6:0] _0048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2603" *)
  wire _0049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2568" *)
  wire [6:0] _0050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2603" *)
  wire _0051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2664" *)
  wire [6:0] _0052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2699" *)
  wire _0053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2664" *)
  wire [6:0] _0054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2699" *)
  wire _0055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2664" *)
  wire [6:0] _0056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2699" *)
  wire _0057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2760" *)
  wire [6:0] _0058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2795" *)
  wire _0059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2760" *)
  wire [6:0] _0060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2795" *)
  wire _0061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2760" *)
  wire [6:0] _0062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2795" *)
  wire _0063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2856" *)
  wire [6:0] _0064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2891" *)
  wire _0065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2856" *)
  wire [6:0] _0066_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2891" *)
  wire _0067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2856" *)
  wire [6:0] _0068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2891" *)
  wire _0069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2952" *)
  wire [6:0] _0070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2987" *)
  wire _0071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2952" *)
  wire [6:0] _0072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2987" *)
  wire _0073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2952" *)
  wire [6:0] _0074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2987" *)
  wire _0075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3048" *)
  wire [6:0] _0076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3083" *)
  wire _0077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3048" *)
  wire [6:0] _0078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3083" *)
  wire _0079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3048" *)
  wire [6:0] _0080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3083" *)
  wire _0081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3144" *)
  wire [6:0] _0082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3179" *)
  wire _0083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3144" *)
  wire [6:0] _0084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3179" *)
  wire _0085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3144" *)
  wire [6:0] _0086_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3179" *)
  wire _0087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3240" *)
  wire [6:0] _0088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3275" *)
  wire _0089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3240" *)
  wire [6:0] _0090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3275" *)
  wire _0091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3240" *)
  wire [6:0] _0092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3275" *)
  wire _0093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3336" *)
  wire [6:0] _0094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3371" *)
  wire _0095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3336" *)
  wire [6:0] _0096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3371" *)
  wire _0097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3336" *)
  wire [6:0] _0098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3371" *)
  wire _0099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3432" *)
  wire [6:0] _0100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3467" *)
  wire _0101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3432" *)
  wire [6:0] _0102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3467" *)
  wire _0103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3432" *)
  wire [6:0] _0104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3467" *)
  wire _0105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2070" *)
  wire [9:0] _0106_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2275" *)
  wire [7:0] _0116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2260" *)
  wire [9:0] _0117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0126_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0146_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0166_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0186_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0203_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0208_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0209_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0210_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0211_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0212_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0213_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0214_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0215_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0216_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0217_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0218_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0232_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0233_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0234_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0235_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0236_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0237_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0238_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0239_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0240_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0241_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0242_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0243_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0244_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0245_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0246_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0247_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0248_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0249_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0250_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0251_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0252_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0253_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0254_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0255_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0256_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0257_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0258_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0259_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0260_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0261_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0262_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0263_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0264_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0265_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0266_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0267_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0268_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0269_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0270_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0271_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0272_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0273_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0274_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0275_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0276_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0277_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0278_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0279_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0280_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0281_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0282_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0283_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0284_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0285_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0286_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0287_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0288_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0289_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0290_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0291_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0292_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0293_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0294_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0295_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0296_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0297_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0298_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0299_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0300_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0301_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0302_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0303_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0304_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0305_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0306_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0307_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0308_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0309_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0310_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0311_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0312_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0313_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0314_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0315_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0316_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0317_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0318_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0319_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0320_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0321_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0322_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0323_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0324_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0325_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0326_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0327_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0328_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0329_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0330_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0331_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0332_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0333_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0334_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0335_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0336_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0337_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0338_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0339_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0340_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0341_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0342_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0343_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0344_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0345_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0346_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0347_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0348_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0349_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0350_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0351_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0352_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0353_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0354_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0355_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0356_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0357_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0358_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0359_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0360_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0361_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0362_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0363_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0364_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0365_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0366_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0367_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0368_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0369_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0370_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0371_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:222" *)
  wire _0372_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:127" *)
  wire [8:0] _0373_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2114" *)
  wire [8:0] _0374_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2117" *)
  wire [8:0] _0375_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2120" *)
  wire [8:0] _0376_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2123" *)
  wire [8:0] _0377_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2126" *)
  wire [8:0] _0378_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2129" *)
  wire [8:0] _0379_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2132" *)
  wire [8:0] _0380_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2135" *)
  wire [8:0] _0381_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2138" *)
  wire [8:0] _0382_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2141" *)
  wire [8:0] _0383_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1001" *)
  wire _0384_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1004" *)
  wire _0385_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1006" *)
  wire _0386_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1009" *)
  wire _0387_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1011" *)
  wire _0388_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1014" *)
  wire _0389_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1016" *)
  wire _0390_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1019" *)
  wire _0391_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1021" *)
  wire _0392_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1024" *)
  wire _0393_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1026" *)
  wire _0394_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1029" *)
  wire _0395_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1031" *)
  wire _0396_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1034" *)
  wire _0397_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1036" *)
  wire _0398_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1039" *)
  wire _0399_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1041" *)
  wire _0400_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1044" *)
  wire _0401_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1046" *)
  wire _0402_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1049" *)
  wire _0403_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1051" *)
  wire _0404_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1054" *)
  wire _0405_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1056" *)
  wire _0406_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1059" *)
  wire _0407_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1061" *)
  wire _0408_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1064" *)
  wire _0409_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1066" *)
  wire _0410_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1069" *)
  wire _0411_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1071" *)
  wire _0412_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1074" *)
  wire _0413_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1076" *)
  wire _0414_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1079" *)
  wire _0415_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1081" *)
  wire _0416_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1084" *)
  wire _0417_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1086" *)
  wire _0418_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1089" *)
  wire _0419_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1091" *)
  wire _0420_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1094" *)
  wire _0421_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1096" *)
  wire _0422_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1099" *)
  wire _0423_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1101" *)
  wire _0424_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1104" *)
  wire _0425_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1106" *)
  wire _0426_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1109" *)
  wire _0427_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1111" *)
  wire _0428_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1114" *)
  wire _0429_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1116" *)
  wire _0430_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1119" *)
  wire _0431_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1121" *)
  wire _0432_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1124" *)
  wire _0433_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1126" *)
  wire _0434_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1129" *)
  wire _0435_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1131" *)
  wire _0436_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1134" *)
  wire _0437_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1136" *)
  wire _0438_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1139" *)
  wire _0439_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1141" *)
  wire _0440_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1144" *)
  wire _0441_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1146" *)
  wire _0442_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1149" *)
  wire _0443_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1151" *)
  wire _0444_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1154" *)
  wire _0445_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1156" *)
  wire _0446_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1159" *)
  wire _0447_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1161" *)
  wire _0448_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1164" *)
  wire _0449_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1166" *)
  wire _0450_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1169" *)
  wire _0451_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1171" *)
  wire _0452_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1174" *)
  wire _0453_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1176" *)
  wire _0454_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1179" *)
  wire _0455_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1181" *)
  wire _0456_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1184" *)
  wire _0457_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1186" *)
  wire _0458_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1189" *)
  wire _0459_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1191" *)
  wire _0460_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1194" *)
  wire _0461_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1196" *)
  wire _0462_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1199" *)
  wire _0463_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1201" *)
  wire _0464_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1204" *)
  wire _0465_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1206" *)
  wire _0466_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1209" *)
  wire _0467_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1211" *)
  wire _0468_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1214" *)
  wire _0469_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1216" *)
  wire _0470_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1219" *)
  wire _0471_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1221" *)
  wire _0472_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1224" *)
  wire _0473_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1226" *)
  wire _0474_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1229" *)
  wire _0475_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1231" *)
  wire _0476_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1234" *)
  wire _0477_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1236" *)
  wire _0478_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1239" *)
  wire _0479_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1241" *)
  wire _0480_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1244" *)
  wire _0481_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1246" *)
  wire _0482_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1249" *)
  wire _0483_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1251" *)
  wire _0484_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1254" *)
  wire _0485_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1256" *)
  wire _0486_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1259" *)
  wire _0487_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1261" *)
  wire _0488_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1264" *)
  wire _0489_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1266" *)
  wire _0490_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1269" *)
  wire _0491_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1271" *)
  wire _0492_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1274" *)
  wire _0493_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1276" *)
  wire _0494_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1279" *)
  wire _0495_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1281" *)
  wire _0496_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1284" *)
  wire _0497_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1286" *)
  wire _0498_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1289" *)
  wire _0499_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1291" *)
  wire _0500_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1294" *)
  wire _0501_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1296" *)
  wire _0502_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1299" *)
  wire _0503_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1301" *)
  wire _0504_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1304" *)
  wire _0505_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1306" *)
  wire _0506_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1309" *)
  wire _0507_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1311" *)
  wire _0508_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1314" *)
  wire _0509_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1316" *)
  wire _0510_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1319" *)
  wire _0511_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1321" *)
  wire _0512_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1324" *)
  wire _0513_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1326" *)
  wire _0514_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1329" *)
  wire _0515_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1331" *)
  wire _0516_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1334" *)
  wire _0517_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1336" *)
  wire _0518_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1339" *)
  wire _0519_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1341" *)
  wire _0520_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1344" *)
  wire _0521_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1346" *)
  wire _0522_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1349" *)
  wire _0523_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1351" *)
  wire _0524_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1354" *)
  wire _0525_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1356" *)
  wire _0526_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1359" *)
  wire _0527_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1361" *)
  wire _0528_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1364" *)
  wire _0529_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1366" *)
  wire _0530_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1369" *)
  wire _0531_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1371" *)
  wire _0532_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1374" *)
  wire _0533_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1376" *)
  wire _0534_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1379" *)
  wire _0535_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1381" *)
  wire _0536_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1384" *)
  wire _0537_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1386" *)
  wire _0538_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1389" *)
  wire _0539_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1391" *)
  wire _0540_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1394" *)
  wire _0541_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1396" *)
  wire _0542_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1399" *)
  wire _0543_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1401" *)
  wire _0544_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1404" *)
  wire _0545_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1406" *)
  wire _0546_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1409" *)
  wire _0547_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1411" *)
  wire _0548_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1414" *)
  wire _0549_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1416" *)
  wire _0550_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1419" *)
  wire _0551_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1421" *)
  wire _0552_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1424" *)
  wire _0553_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1426" *)
  wire _0554_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1429" *)
  wire _0555_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1431" *)
  wire _0556_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1434" *)
  wire _0557_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1436" *)
  wire _0558_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1439" *)
  wire _0559_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1441" *)
  wire _0560_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1444" *)
  wire _0561_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1446" *)
  wire _0562_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1449" *)
  wire _0563_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1451" *)
  wire _0564_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1454" *)
  wire _0565_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1456" *)
  wire _0566_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1459" *)
  wire _0567_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1461" *)
  wire _0568_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1464" *)
  wire _0569_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1466" *)
  wire _0570_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1469" *)
  wire _0571_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1471" *)
  wire _0572_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1474" *)
  wire _0573_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1476" *)
  wire _0574_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1479" *)
  wire _0575_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1481" *)
  wire _0576_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1484" *)
  wire _0577_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1486" *)
  wire _0578_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1489" *)
  wire _0579_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1491" *)
  wire _0580_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1494" *)
  wire _0581_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1496" *)
  wire _0582_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2013" *)
  wire _0583_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2014" *)
  wire _0584_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2015" *)
  wire _0585_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2016" *)
  wire _0586_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2017" *)
  wire _0587_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2018" *)
  wire _0588_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2019" *)
  wire _0589_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2020" *)
  wire _0590_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2021" *)
  wire _0591_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2022" *)
  wire _0592_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2037" *)
  wire _0593_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2038" *)
  wire _0594_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2039" *)
  wire _0595_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2040" *)
  wire _0596_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2041" *)
  wire _0597_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2042" *)
  wire _0598_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2043" *)
  wire _0599_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2044" *)
  wire _0600_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2045" *)
  wire _0601_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2046" *)
  wire _0602_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:224" *)
  wire _0603_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:226" *)
  wire _0604_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2285" *)
  wire _0605_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *)
  wire _0606_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:229" *)
  wire _0607_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2300" *)
  wire _0608_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *)
  wire _0609_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:231" *)
  wire _0610_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2315" *)
  wire _0611_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *)
  wire _0612_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2330" *)
  wire _0613_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *)
  wire _0614_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:234" *)
  wire _0615_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2345" *)
  wire _0616_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *)
  wire _0617_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:236" *)
  wire _0618_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2360" *)
  wire _0619_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *)
  wire _0620_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2375" *)
  wire _0621_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *)
  wire _0622_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:239" *)
  wire _0623_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2390" *)
  wire _0624_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *)
  wire _0625_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2405" *)
  wire _0626_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *)
  wire _0627_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:241" *)
  wire _0628_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2420" *)
  wire _0629_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *)
  wire _0630_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:244" *)
  wire _0631_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:246" *)
  wire _0632_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:249" *)
  wire _0633_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:251" *)
  wire _0634_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:254" *)
  wire _0635_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:256" *)
  wire _0636_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:259" *)
  wire _0637_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:261" *)
  wire _0638_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _0639_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:264" *)
  wire _0640_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:266" *)
  wire _0641_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:269" *)
  wire _0642_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:271" *)
  wire _0643_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _0644_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:274" *)
  wire _0645_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:276" *)
  wire _0646_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:279" *)
  wire _0647_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:281" *)
  wire _0648_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _0649_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:284" *)
  wire _0650_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:286" *)
  wire _0651_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:289" *)
  wire _0652_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:291" *)
  wire _0653_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _0654_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:294" *)
  wire _0655_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:296" *)
  wire _0656_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:299" *)
  wire _0657_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:301" *)
  wire _0658_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _0659_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:304" *)
  wire _0660_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:306" *)
  wire _0661_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:309" *)
  wire _0662_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _0663_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:311" *)
  wire _0664_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:314" *)
  wire _0665_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:316" *)
  wire _0666_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:319" *)
  wire _0667_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _0668_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:321" *)
  wire _0669_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:324" *)
  wire _0670_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:326" *)
  wire _0671_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:329" *)
  wire _0672_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _0673_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:331" *)
  wire _0674_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:334" *)
  wire _0675_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:336" *)
  wire _0676_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:339" *)
  wire _0677_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _0678_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:341" *)
  wire _0679_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:344" *)
  wire _0680_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:346" *)
  wire _0681_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:349" *)
  wire _0682_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _0683_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:351" *)
  wire _0684_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *)
  wire _0685_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *)
  wire _0686_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *)
  wire _0687_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _0688_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _0689_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _0690_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _0691_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _0692_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _0693_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3522" *)
  wire _0694_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:354" *)
  wire _0695_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:356" *)
  wire _0696_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:359" *)
  wire _0697_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:361" *)
  wire _0698_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:364" *)
  wire _0699_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:366" *)
  wire _0700_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:369" *)
  wire _0701_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:371" *)
  wire _0702_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:374" *)
  wire _0703_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:376" *)
  wire _0704_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:379" *)
  wire _0705_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:381" *)
  wire _0706_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:384" *)
  wire _0707_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:386" *)
  wire _0708_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:389" *)
  wire _0709_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:391" *)
  wire _0710_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:394" *)
  wire _0711_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:396" *)
  wire _0712_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:399" *)
  wire _0713_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:401" *)
  wire _0714_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:404" *)
  wire _0715_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:406" *)
  wire _0716_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:409" *)
  wire _0717_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:411" *)
  wire _0718_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:414" *)
  wire _0719_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:416" *)
  wire _0720_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:419" *)
  wire _0721_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:421" *)
  wire _0722_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:424" *)
  wire _0723_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:426" *)
  wire _0724_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:429" *)
  wire _0725_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:431" *)
  wire _0726_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:434" *)
  wire _0727_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:436" *)
  wire _0728_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:439" *)
  wire _0729_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:441" *)
  wire _0730_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:444" *)
  wire _0731_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:446" *)
  wire _0732_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:449" *)
  wire _0733_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:451" *)
  wire _0734_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:454" *)
  wire _0735_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:456" *)
  wire _0736_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:459" *)
  wire _0737_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:461" *)
  wire _0738_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:464" *)
  wire _0739_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:466" *)
  wire _0740_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:469" *)
  wire _0741_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:471" *)
  wire _0742_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:474" *)
  wire _0743_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:476" *)
  wire _0744_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:479" *)
  wire _0745_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:481" *)
  wire _0746_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:484" *)
  wire _0747_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:486" *)
  wire _0748_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:489" *)
  wire _0749_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:491" *)
  wire _0750_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:494" *)
  wire _0751_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:496" *)
  wire _0752_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:499" *)
  wire _0753_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:501" *)
  wire _0754_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:504" *)
  wire _0755_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:506" *)
  wire _0756_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:509" *)
  wire _0757_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:511" *)
  wire _0758_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:514" *)
  wire _0759_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:516" *)
  wire _0760_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:519" *)
  wire _0761_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:521" *)
  wire _0762_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:524" *)
  wire _0763_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:526" *)
  wire _0764_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:529" *)
  wire _0765_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:531" *)
  wire _0766_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:534" *)
  wire _0767_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:536" *)
  wire _0768_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:539" *)
  wire _0769_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:541" *)
  wire _0770_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:544" *)
  wire _0771_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:546" *)
  wire _0772_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:549" *)
  wire _0773_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:551" *)
  wire _0774_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:554" *)
  wire _0775_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:556" *)
  wire _0776_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:559" *)
  wire _0777_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:561" *)
  wire _0778_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:564" *)
  wire _0779_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:566" *)
  wire _0780_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:569" *)
  wire _0781_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:571" *)
  wire _0782_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:574" *)
  wire _0783_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:576" *)
  wire _0784_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:579" *)
  wire _0785_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:581" *)
  wire _0786_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:584" *)
  wire _0787_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:586" *)
  wire _0788_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:589" *)
  wire _0789_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:591" *)
  wire _0790_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:594" *)
  wire _0791_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:596" *)
  wire _0792_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:599" *)
  wire _0793_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:601" *)
  wire _0794_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:604" *)
  wire _0795_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:606" *)
  wire _0796_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:609" *)
  wire _0797_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:611" *)
  wire _0798_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:614" *)
  wire _0799_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:616" *)
  wire _0800_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:619" *)
  wire _0801_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:621" *)
  wire _0802_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:624" *)
  wire _0803_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:626" *)
  wire _0804_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:629" *)
  wire _0805_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:631" *)
  wire _0806_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:634" *)
  wire _0807_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:636" *)
  wire _0808_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:639" *)
  wire _0809_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:641" *)
  wire _0810_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:644" *)
  wire _0811_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:646" *)
  wire _0812_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:649" *)
  wire _0813_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:651" *)
  wire _0814_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:654" *)
  wire _0815_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:656" *)
  wire _0816_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:659" *)
  wire _0817_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:661" *)
  wire _0818_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:664" *)
  wire _0819_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:666" *)
  wire _0820_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:669" *)
  wire _0821_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:671" *)
  wire _0822_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:674" *)
  wire _0823_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:676" *)
  wire _0824_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:679" *)
  wire _0825_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:681" *)
  wire _0826_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:684" *)
  wire _0827_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:686" *)
  wire _0828_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:689" *)
  wire _0829_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:691" *)
  wire _0830_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:694" *)
  wire _0831_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:696" *)
  wire _0832_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:699" *)
  wire _0833_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:701" *)
  wire _0834_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:704" *)
  wire _0835_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:706" *)
  wire _0836_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:709" *)
  wire _0837_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:711" *)
  wire _0838_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:714" *)
  wire _0839_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:716" *)
  wire _0840_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:719" *)
  wire _0841_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:721" *)
  wire _0842_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:724" *)
  wire _0843_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:726" *)
  wire _0844_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:729" *)
  wire _0845_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:731" *)
  wire _0846_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:734" *)
  wire _0847_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:736" *)
  wire _0848_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:739" *)
  wire _0849_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:741" *)
  wire _0850_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:744" *)
  wire _0851_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:746" *)
  wire _0852_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:749" *)
  wire _0853_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:751" *)
  wire _0854_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:754" *)
  wire _0855_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:756" *)
  wire _0856_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:759" *)
  wire _0857_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:761" *)
  wire _0858_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:764" *)
  wire _0859_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:766" *)
  wire _0860_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:769" *)
  wire _0861_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:771" *)
  wire _0862_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:774" *)
  wire _0863_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:776" *)
  wire _0864_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:779" *)
  wire _0865_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:781" *)
  wire _0866_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:784" *)
  wire _0867_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:786" *)
  wire _0868_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:789" *)
  wire _0869_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:791" *)
  wire _0870_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:794" *)
  wire _0871_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:796" *)
  wire _0872_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:799" *)
  wire _0873_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:801" *)
  wire _0874_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:804" *)
  wire _0875_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:806" *)
  wire _0876_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:809" *)
  wire _0877_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:811" *)
  wire _0878_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:814" *)
  wire _0879_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:816" *)
  wire _0880_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:819" *)
  wire _0881_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:821" *)
  wire _0882_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:824" *)
  wire _0883_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:826" *)
  wire _0884_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:829" *)
  wire _0885_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:831" *)
  wire _0886_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:834" *)
  wire _0887_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:836" *)
  wire _0888_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:839" *)
  wire _0889_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:841" *)
  wire _0890_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:844" *)
  wire _0891_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:846" *)
  wire _0892_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:849" *)
  wire _0893_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:851" *)
  wire _0894_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:854" *)
  wire _0895_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:856" *)
  wire _0896_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:859" *)
  wire _0897_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:861" *)
  wire _0898_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:864" *)
  wire _0899_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:866" *)
  wire _0900_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:869" *)
  wire _0901_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:871" *)
  wire _0902_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:874" *)
  wire _0903_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:876" *)
  wire _0904_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:879" *)
  wire _0905_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:881" *)
  wire _0906_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:884" *)
  wire _0907_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:886" *)
  wire _0908_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:889" *)
  wire _0909_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:891" *)
  wire _0910_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:894" *)
  wire _0911_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:896" *)
  wire _0912_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:899" *)
  wire _0913_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:901" *)
  wire _0914_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:904" *)
  wire _0915_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:906" *)
  wire _0916_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:909" *)
  wire _0917_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:911" *)
  wire _0918_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:914" *)
  wire _0919_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:916" *)
  wire _0920_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:919" *)
  wire _0921_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:921" *)
  wire _0922_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:924" *)
  wire _0923_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:926" *)
  wire _0924_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:929" *)
  wire _0925_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:931" *)
  wire _0926_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:934" *)
  wire _0927_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:936" *)
  wire _0928_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:939" *)
  wire _0929_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:941" *)
  wire _0930_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:944" *)
  wire _0931_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:946" *)
  wire _0932_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:949" *)
  wire _0933_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:951" *)
  wire _0934_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:954" *)
  wire _0935_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:956" *)
  wire _0936_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:959" *)
  wire _0937_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:961" *)
  wire _0938_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:964" *)
  wire _0939_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:966" *)
  wire _0940_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:969" *)
  wire _0941_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:971" *)
  wire _0942_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:974" *)
  wire _0943_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:976" *)
  wire _0944_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:979" *)
  wire _0945_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:981" *)
  wire _0946_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:984" *)
  wire _0947_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:986" *)
  wire _0948_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:989" *)
  wire _0949_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:991" *)
  wire _0950_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:994" *)
  wire _0951_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:996" *)
  wire _0952_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:999" *)
  wire _0953_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2250" *)
  wire _0954_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2251" *)
  wire _0955_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2252" *)
  wire _0956_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2253" *)
  wire _0957_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2254" *)
  wire _0958_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2255" *)
  wire _0959_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2256" *)
  wire _0960_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2257" *)
  wire _0961_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2258" *)
  wire _0962_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2259" *)
  wire _0963_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1001" *)
  wire _0964_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1004" *)
  wire _0965_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1006" *)
  wire _0966_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1009" *)
  wire _0967_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1011" *)
  wire _0968_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1014" *)
  wire _0969_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1016" *)
  wire _0970_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1019" *)
  wire _0971_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1021" *)
  wire _0972_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1024" *)
  wire _0973_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1026" *)
  wire _0974_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1029" *)
  wire _0975_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1031" *)
  wire _0976_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1034" *)
  wire _0977_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1036" *)
  wire _0978_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1039" *)
  wire _0979_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1041" *)
  wire _0980_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1044" *)
  wire _0981_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1046" *)
  wire _0982_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1049" *)
  wire _0983_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1051" *)
  wire _0984_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1054" *)
  wire _0985_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1056" *)
  wire _0986_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1059" *)
  wire _0987_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1061" *)
  wire _0988_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1064" *)
  wire _0989_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1066" *)
  wire _0990_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1069" *)
  wire _0991_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1071" *)
  wire _0992_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1074" *)
  wire _0993_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1076" *)
  wire _0994_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1079" *)
  wire _0995_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1081" *)
  wire _0996_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1084" *)
  wire _0997_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1086" *)
  wire _0998_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1089" *)
  wire _0999_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1091" *)
  wire _1000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1094" *)
  wire _1001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1096" *)
  wire _1002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1099" *)
  wire _1003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1101" *)
  wire _1004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1104" *)
  wire _1005_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1106" *)
  wire _1006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1109" *)
  wire _1007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1111" *)
  wire _1008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1114" *)
  wire _1009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1116" *)
  wire _1010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1119" *)
  wire _1011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1121" *)
  wire _1012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1124" *)
  wire _1013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1126" *)
  wire _1014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1129" *)
  wire _1015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1131" *)
  wire _1016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1134" *)
  wire _1017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1136" *)
  wire _1018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1139" *)
  wire _1019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1141" *)
  wire _1020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1144" *)
  wire _1021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1146" *)
  wire _1022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1149" *)
  wire _1023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1151" *)
  wire _1024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1154" *)
  wire _1025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1156" *)
  wire _1026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1159" *)
  wire _1027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1161" *)
  wire _1028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1164" *)
  wire _1029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1166" *)
  wire _1030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1169" *)
  wire _1031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1171" *)
  wire _1032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1174" *)
  wire _1033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1176" *)
  wire _1034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1179" *)
  wire _1035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1181" *)
  wire _1036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1184" *)
  wire _1037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1186" *)
  wire _1038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1189" *)
  wire _1039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1191" *)
  wire _1040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1194" *)
  wire _1041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1196" *)
  wire _1042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1199" *)
  wire _1043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1201" *)
  wire _1044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1204" *)
  wire _1045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1206" *)
  wire _1046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1209" *)
  wire _1047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1211" *)
  wire _1048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1214" *)
  wire _1049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1216" *)
  wire _1050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1219" *)
  wire _1051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1221" *)
  wire _1052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1224" *)
  wire _1053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1226" *)
  wire _1054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1229" *)
  wire _1055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1231" *)
  wire _1056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1234" *)
  wire _1057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1236" *)
  wire _1058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1239" *)
  wire _1059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1241" *)
  wire _1060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1244" *)
  wire _1061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1246" *)
  wire _1062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1249" *)
  wire _1063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1251" *)
  wire _1064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1254" *)
  wire _1065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1256" *)
  wire _1066_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1259" *)
  wire _1067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1261" *)
  wire _1068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1264" *)
  wire _1069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1266" *)
  wire _1070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1269" *)
  wire _1071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1271" *)
  wire _1072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1274" *)
  wire _1073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1276" *)
  wire _1074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1279" *)
  wire _1075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1281" *)
  wire _1076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1284" *)
  wire _1077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1286" *)
  wire _1078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1289" *)
  wire _1079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1291" *)
  wire _1080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1294" *)
  wire _1081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1296" *)
  wire _1082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1299" *)
  wire _1083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1301" *)
  wire _1084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1304" *)
  wire _1085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1306" *)
  wire _1086_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1309" *)
  wire _1087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1311" *)
  wire _1088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1314" *)
  wire _1089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1316" *)
  wire _1090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1319" *)
  wire _1091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1321" *)
  wire _1092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1324" *)
  wire _1093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1326" *)
  wire _1094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1329" *)
  wire _1095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1331" *)
  wire _1096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1334" *)
  wire _1097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1336" *)
  wire _1098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1339" *)
  wire _1099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1341" *)
  wire _1100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1344" *)
  wire _1101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1346" *)
  wire _1102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1349" *)
  wire _1103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1351" *)
  wire _1104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1354" *)
  wire _1105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1356" *)
  wire _1106_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1359" *)
  wire _1107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1361" *)
  wire _1108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1364" *)
  wire _1109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1366" *)
  wire _1110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1369" *)
  wire _1111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1371" *)
  wire _1112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1374" *)
  wire _1113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1376" *)
  wire _1114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1379" *)
  wire _1115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1381" *)
  wire _1116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1384" *)
  wire _1117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1386" *)
  wire _1118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1389" *)
  wire _1119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1391" *)
  wire _1120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1394" *)
  wire _1121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1396" *)
  wire _1122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1399" *)
  wire _1123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1401" *)
  wire _1124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1404" *)
  wire _1125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1406" *)
  wire _1126_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1409" *)
  wire _1127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1411" *)
  wire _1128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1414" *)
  wire _1129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1416" *)
  wire _1130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1419" *)
  wire _1131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1421" *)
  wire _1132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1424" *)
  wire _1133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1426" *)
  wire _1134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1429" *)
  wire _1135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1431" *)
  wire _1136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1434" *)
  wire _1137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1436" *)
  wire _1138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1439" *)
  wire _1139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1441" *)
  wire _1140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1444" *)
  wire _1141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1446" *)
  wire _1142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1449" *)
  wire _1143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1451" *)
  wire _1144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1454" *)
  wire _1145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1456" *)
  wire _1146_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1459" *)
  wire _1147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1461" *)
  wire _1148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1464" *)
  wire _1149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1466" *)
  wire _1150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1469" *)
  wire _1151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1471" *)
  wire _1152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1474" *)
  wire _1153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1476" *)
  wire _1154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1479" *)
  wire _1155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1481" *)
  wire _1156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1484" *)
  wire _1157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1486" *)
  wire _1158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1489" *)
  wire _1159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1491" *)
  wire _1160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1494" *)
  wire _1161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1496" *)
  wire _1162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:224" *)
  wire _1163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:226" *)
  wire _1164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2285" *)
  wire _1165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *)
  wire _1166_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *)
  wire _1167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:229" *)
  wire _1168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2300" *)
  wire _1169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *)
  wire _1170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *)
  wire _1171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:231" *)
  wire _1172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2315" *)
  wire _1173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *)
  wire _1174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *)
  wire _1175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2330" *)
  wire _1176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *)
  wire _1177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *)
  wire _1178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:234" *)
  wire _1179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2345" *)
  wire _1180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *)
  wire _1181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *)
  wire _1182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:236" *)
  wire _1183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2360" *)
  wire _1184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *)
  wire _1185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *)
  wire _1186_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2375" *)
  wire _1187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *)
  wire _1188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *)
  wire _1189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:239" *)
  wire _1190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2390" *)
  wire _1191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *)
  wire _1192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *)
  wire _1193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2405" *)
  wire _1194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *)
  wire _1195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *)
  wire _1196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:241" *)
  wire _1197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2420" *)
  wire _1198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *)
  wire _1199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *)
  wire _1200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:244" *)
  wire _1201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2457" *)
  wire _1202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2458" *)
  wire _1203_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2459" *)
  wire _1204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:246" *)
  wire _1205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2460" *)
  wire _1206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2461" *)
  wire _1207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2462" *)
  wire _1208_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2463" *)
  wire _1209_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2464" *)
  wire _1210_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2465" *)
  wire _1211_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2466" *)
  wire _1212_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2474" *)
  wire _1213_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2475" *)
  wire _1214_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2476" *)
  wire _1215_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2477" *)
  wire _1216_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2478" *)
  wire _1217_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2479" *)
  wire _1218_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2480" *)
  wire _1219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2481" *)
  wire _1220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2482" *)
  wire _1221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2483" *)
  wire _1222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:249" *)
  wire _1223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2491" *)
  wire _1224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2492" *)
  wire _1225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2493" *)
  wire _1226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2494" *)
  wire _1227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2495" *)
  wire _1228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2496" *)
  wire _1229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2497" *)
  wire _1230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2498" *)
  wire _1231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2499" *)
  wire _1232_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2500" *)
  wire _1233_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:251" *)
  wire _1234_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:254" *)
  wire _1235_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:256" *)
  wire _1236_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _1237_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _1238_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _1239_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2571" *)
  wire _1240_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *)
  wire _1241_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *)
  wire _1242_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2583" *)
  wire _1243_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:259" *)
  wire _1244_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *)
  wire _1245_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *)
  wire _1246_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *)
  wire _1247_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *)
  wire _1248_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:261" *)
  wire _1249_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *)
  wire _1250_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2612" *)
  wire _1251_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _1252_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _1253_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _1254_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _1255_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _1256_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _1257_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _1258_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:264" *)
  wire _1259_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:266" *)
  wire _1260_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _1261_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _1262_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _1263_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2667" *)
  wire _1264_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *)
  wire _1265_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *)
  wire _1266_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2679" *)
  wire _1267_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *)
  wire _1268_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *)
  wire _1269_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *)
  wire _1270_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:269" *)
  wire _1271_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *)
  wire _1272_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *)
  wire _1273_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2708" *)
  wire _1274_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:271" *)
  wire _1275_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _1276_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _1277_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _1278_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _1279_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _1280_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _1281_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _1282_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:274" *)
  wire _1283_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:276" *)
  wire _1284_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _1285_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _1286_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _1287_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2763" *)
  wire _1288_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *)
  wire _1289_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *)
  wire _1290_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2775" *)
  wire _1291_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *)
  wire _1292_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *)
  wire _1293_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *)
  wire _1294_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:279" *)
  wire _1295_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *)
  wire _1296_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *)
  wire _1297_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2804" *)
  wire _1298_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:281" *)
  wire _1299_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _1300_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _1301_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _1302_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _1303_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _1304_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _1305_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _1306_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:284" *)
  wire _1307_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _1308_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _1309_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _1310_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2859" *)
  wire _1311_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:286" *)
  wire _1312_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *)
  wire _1313_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *)
  wire _1314_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2871" *)
  wire _1315_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *)
  wire _1316_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *)
  wire _1317_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *)
  wire _1318_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:289" *)
  wire _1319_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *)
  wire _1320_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *)
  wire _1321_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2900" *)
  wire _1322_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:291" *)
  wire _1323_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _1324_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _1325_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _1326_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _1327_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _1328_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _1329_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _1330_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:294" *)
  wire _1331_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _1332_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _1333_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _1334_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2955" *)
  wire _1335_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:296" *)
  wire _1336_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *)
  wire _1337_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *)
  wire _1338_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2967" *)
  wire _1339_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *)
  wire _1340_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *)
  wire _1341_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *)
  wire _1342_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:299" *)
  wire _1343_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *)
  wire _1344_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *)
  wire _1345_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2996" *)
  wire _1346_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _1347_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:301" *)
  wire _1348_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _1349_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _1350_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _1351_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _1352_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _1353_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _1354_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:304" *)
  wire _1355_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _1356_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _1357_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _1358_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3051" *)
  wire _1359_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:306" *)
  wire _1360_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *)
  wire _1361_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *)
  wire _1362_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3063" *)
  wire _1363_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *)
  wire _1364_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *)
  wire _1365_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *)
  wire _1366_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *)
  wire _1367_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:309" *)
  wire _1368_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *)
  wire _1369_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3092" *)
  wire _1370_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _1371_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _1372_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _1373_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _1374_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _1375_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _1376_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _1377_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:311" *)
  wire _1378_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:314" *)
  wire _1379_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _1380_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _1381_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _1382_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3147" *)
  wire _1383_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *)
  wire _1384_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *)
  wire _1385_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3159" *)
  wire _1386_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:316" *)
  wire _1387_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *)
  wire _1388_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *)
  wire _1389_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *)
  wire _1390_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *)
  wire _1391_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *)
  wire _1392_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3188" *)
  wire _1393_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:319" *)
  wire _1394_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _1395_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _1396_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _1397_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _1398_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _1399_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _1400_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _1401_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:321" *)
  wire _1402_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:324" *)
  wire _1403_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _1404_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _1405_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _1406_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3243" *)
  wire _1407_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *)
  wire _1408_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *)
  wire _1409_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3255" *)
  wire _1410_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:326" *)
  wire _1411_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *)
  wire _1412_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *)
  wire _1413_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *)
  wire _1414_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *)
  wire _1415_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *)
  wire _1416_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3284" *)
  wire _1417_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:329" *)
  wire _1418_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _1419_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _1420_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _1421_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _1422_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _1423_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _1424_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _1425_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:331" *)
  wire _1426_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _1427_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _1428_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _1429_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3339" *)
  wire _1430_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:334" *)
  wire _1431_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *)
  wire _1432_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *)
  wire _1433_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3351" *)
  wire _1434_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:336" *)
  wire _1435_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *)
  wire _1436_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *)
  wire _1437_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *)
  wire _1438_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *)
  wire _1439_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *)
  wire _1440_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3380" *)
  wire _1441_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:339" *)
  wire _1442_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _1443_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _1444_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _1445_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _1446_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _1447_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _1448_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _1449_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:341" *)
  wire _1450_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _1451_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _1452_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _1453_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3435" *)
  wire _1454_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:344" *)
  wire _1455_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *)
  wire _1456_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *)
  wire _1457_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3447" *)
  wire _1458_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *)
  wire _1459_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *)
  wire _1460_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *)
  wire _1461_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:346" *)
  wire _1462_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *)
  wire _1463_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *)
  wire _1464_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3476" *)
  wire _1465_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _1466_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:349" *)
  wire _1467_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _1468_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _1469_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _1470_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _1471_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _1472_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _1473_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:351" *)
  wire _1474_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *)
  wire _1475_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *)
  wire _1476_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *)
  wire _1477_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *)
  wire _1478_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *)
  wire _1479_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *)
  wire _1480_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _1481_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _1482_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _1483_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _1484_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _1485_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _1486_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _1487_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _1488_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _1489_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1490_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1491_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1492_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1493_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1494_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _1495_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1496_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1497_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1498_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1499_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1500_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1501_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _1502_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1503_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1504_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1505_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1506_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1507_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1508_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1509_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _1510_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1511_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1512_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1513_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1514_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1515_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1516_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1517_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1518_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _1519_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *)
  wire _1520_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *)
  wire _1521_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *)
  wire _1522_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *)
  wire _1523_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *)
  wire _1524_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *)
  wire _1525_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *)
  wire _1526_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *)
  wire _1527_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *)
  wire _1528_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *)
  wire _1529_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *)
  wire _1530_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *)
  wire _1531_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *)
  wire _1532_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *)
  wire _1533_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1534_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1535_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1536_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1537_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1538_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *)
  wire _1539_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1540_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1541_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1542_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1543_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1544_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1545_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *)
  wire _1546_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1547_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1548_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1549_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1550_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1551_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1552_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1553_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *)
  wire _1554_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1555_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1556_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1557_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1558_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1559_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1560_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1561_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1562_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *)
  wire _1563_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3533" *)
  wire _1564_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *)
  wire _1565_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *)
  wire _1566_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *)
  wire _1567_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *)
  wire _1568_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *)
  wire _1569_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *)
  wire _1570_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *)
  wire _1571_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *)
  wire _1572_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *)
  wire _1573_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *)
  wire _1574_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *)
  wire _1575_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *)
  wire _1576_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1577_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1578_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1579_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1580_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1581_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *)
  wire _1582_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1583_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1584_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1585_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1586_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1587_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1588_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *)
  wire _1589_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:354" *)
  wire _1590_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1591_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1592_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1593_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1594_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1595_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1596_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1597_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *)
  wire _1598_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1599_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1600_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1601_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1602_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1603_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1604_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1605_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1606_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *)
  wire _1607_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3543" *)
  wire _1608_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3544" *)
  wire _1609_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3544" *)
  wire _1610_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *)
  wire _1611_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *)
  wire _1612_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *)
  wire _1613_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *)
  wire _1614_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *)
  wire _1615_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *)
  wire _1616_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *)
  wire _1617_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *)
  wire _1618_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *)
  wire _1619_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1620_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1621_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1622_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1623_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1624_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *)
  wire _1625_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1626_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1627_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1628_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1629_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1630_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1631_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *)
  wire _1632_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1633_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1634_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1635_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1636_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1637_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1638_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1639_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *)
  wire _1640_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1641_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1642_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1643_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1644_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1645_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1646_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1647_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1648_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *)
  wire _1649_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3553" *)
  wire _1650_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3554" *)
  wire _1651_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3554" *)
  wire _1652_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *)
  wire _1653_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *)
  wire _1654_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *)
  wire _1655_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *)
  wire _1656_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *)
  wire _1657_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *)
  wire _1658_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *)
  wire _1659_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *)
  wire _1660_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1661_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1662_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1663_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1664_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1665_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *)
  wire _1666_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1667_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1668_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1669_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1670_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1671_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1672_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *)
  wire _1673_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:356" *)
  wire _1674_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1675_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1676_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1677_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1678_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1679_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1680_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1681_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *)
  wire _1682_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1683_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1684_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1685_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1686_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1687_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1688_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1689_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1690_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *)
  wire _1691_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3563" *)
  wire _1692_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3564" *)
  wire _1693_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3564" *)
  wire _1694_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *)
  wire _1695_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *)
  wire _1696_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *)
  wire _1697_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *)
  wire _1698_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *)
  wire _1699_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *)
  wire _1700_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *)
  wire _1701_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1702_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1703_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1704_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1705_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1706_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *)
  wire _1707_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1708_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1709_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1710_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1711_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1712_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1713_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *)
  wire _1714_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1715_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1716_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1717_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1718_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1719_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1720_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1721_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *)
  wire _1722_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1723_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1724_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1725_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1726_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1727_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1728_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1729_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1730_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *)
  wire _1731_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3573" *)
  wire _1732_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3574" *)
  wire _1733_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3574" *)
  wire _1734_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *)
  wire _1735_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *)
  wire _1736_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *)
  wire _1737_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *)
  wire _1738_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *)
  wire _1739_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *)
  wire _1740_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *)
  wire _1741_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *)
  wire _1742_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *)
  wire _1743_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *)
  wire _1744_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *)
  wire _1745_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *)
  wire _1746_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1747_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1748_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1749_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1750_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1751_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1752_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *)
  wire _1753_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1754_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1755_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1756_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1757_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1758_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1759_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1760_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *)
  wire _1761_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1762_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1763_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1764_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1765_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1766_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1767_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1768_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1769_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *)
  wire _1770_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3583" *)
  wire _1771_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3584" *)
  wire _1772_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3584" *)
  wire _1773_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *)
  wire _1774_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *)
  wire _1775_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *)
  wire _1776_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *)
  wire _1777_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *)
  wire _1778_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *)
  wire _1779_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *)
  wire _1780_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *)
  wire _1781_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *)
  wire _1782_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *)
  wire _1783_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *)
  wire _1784_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *)
  wire _1785_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1786_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1787_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1788_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1789_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1790_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *)
  wire _1791_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:359" *)
  wire _1792_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1793_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1794_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1795_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1796_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1797_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1798_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1799_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *)
  wire _1800_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1801_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1802_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1803_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1804_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1805_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1806_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1807_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1808_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *)
  wire _1809_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3593" *)
  wire _1810_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3594" *)
  wire _1811_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3594" *)
  wire _1812_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *)
  wire _1813_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *)
  wire _1814_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *)
  wire _1815_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *)
  wire _1816_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *)
  wire _1817_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *)
  wire _1818_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *)
  wire _1819_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *)
  wire _1820_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *)
  wire _1821_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *)
  wire _1822_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *)
  wire _1823_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *)
  wire _1824_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1825_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1826_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1827_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1828_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1829_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *)
  wire _1830_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1831_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1832_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1833_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1834_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1835_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1836_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *)
  wire _1837_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1838_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1839_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1840_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1841_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1842_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1843_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1844_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1845_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *)
  wire _1846_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3603" *)
  wire _1847_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3604" *)
  wire _1848_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3604" *)
  wire _1849_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *)
  wire _1850_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *)
  wire _1851_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *)
  wire _1852_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *)
  wire _1853_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *)
  wire _1854_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *)
  wire _1855_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *)
  wire _1856_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *)
  wire _1857_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *)
  wire _1858_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *)
  wire _1859_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *)
  wire _1860_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *)
  wire _1861_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1862_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1863_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1864_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1865_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1866_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *)
  wire _1867_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1868_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1869_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1870_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1871_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1872_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1873_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *)
  wire _1874_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:361" *)
  wire _1875_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1876_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1877_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1878_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1879_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1880_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1881_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1882_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *)
  wire _1883_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:364" *)
  wire _1884_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:366" *)
  wire _1885_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:369" *)
  wire _1886_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:371" *)
  wire _1887_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:374" *)
  wire _1888_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:376" *)
  wire _1889_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:379" *)
  wire _1890_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:381" *)
  wire _1891_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:384" *)
  wire _1892_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:386" *)
  wire _1893_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:389" *)
  wire _1894_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:391" *)
  wire _1895_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:394" *)
  wire _1896_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:396" *)
  wire _1897_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:399" *)
  wire _1898_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:401" *)
  wire _1899_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:404" *)
  wire _1900_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:406" *)
  wire _1901_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:409" *)
  wire _1902_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:411" *)
  wire _1903_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:414" *)
  wire _1904_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:416" *)
  wire _1905_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:419" *)
  wire _1906_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:421" *)
  wire _1907_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:424" *)
  wire _1908_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:426" *)
  wire _1909_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:429" *)
  wire _1910_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:431" *)
  wire _1911_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:434" *)
  wire _1912_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:436" *)
  wire _1913_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:439" *)
  wire _1914_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:441" *)
  wire _1915_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:444" *)
  wire _1916_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:446" *)
  wire _1917_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:449" *)
  wire _1918_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:451" *)
  wire _1919_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:454" *)
  wire _1920_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:456" *)
  wire _1921_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:459" *)
  wire _1922_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:461" *)
  wire _1923_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:464" *)
  wire _1924_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:466" *)
  wire _1925_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:469" *)
  wire _1926_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:471" *)
  wire _1927_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:474" *)
  wire _1928_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:476" *)
  wire _1929_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:479" *)
  wire _1930_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:481" *)
  wire _1931_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:484" *)
  wire _1932_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:486" *)
  wire _1933_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:489" *)
  wire _1934_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:491" *)
  wire _1935_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:494" *)
  wire _1936_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:496" *)
  wire _1937_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:499" *)
  wire _1938_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:501" *)
  wire _1939_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:504" *)
  wire _1940_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:506" *)
  wire _1941_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:509" *)
  wire _1942_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:511" *)
  wire _1943_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:514" *)
  wire _1944_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:516" *)
  wire _1945_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:519" *)
  wire _1946_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:521" *)
  wire _1947_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:524" *)
  wire _1948_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:526" *)
  wire _1949_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:529" *)
  wire _1950_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:531" *)
  wire _1951_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:534" *)
  wire _1952_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:536" *)
  wire _1953_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:539" *)
  wire _1954_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:541" *)
  wire _1955_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:544" *)
  wire _1956_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:546" *)
  wire _1957_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:549" *)
  wire _1958_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:551" *)
  wire _1959_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:554" *)
  wire _1960_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:556" *)
  wire _1961_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:559" *)
  wire _1962_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:561" *)
  wire _1963_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:564" *)
  wire _1964_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:566" *)
  wire _1965_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:569" *)
  wire _1966_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:571" *)
  wire _1967_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:574" *)
  wire _1968_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:576" *)
  wire _1969_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:579" *)
  wire _1970_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:581" *)
  wire _1971_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:584" *)
  wire _1972_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:586" *)
  wire _1973_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:589" *)
  wire _1974_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:591" *)
  wire _1975_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:594" *)
  wire _1976_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:596" *)
  wire _1977_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:599" *)
  wire _1978_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:601" *)
  wire _1979_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:604" *)
  wire _1980_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:606" *)
  wire _1981_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:609" *)
  wire _1982_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:611" *)
  wire _1983_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:614" *)
  wire _1984_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:616" *)
  wire _1985_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:619" *)
  wire _1986_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:621" *)
  wire _1987_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:624" *)
  wire _1988_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:626" *)
  wire _1989_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:629" *)
  wire _1990_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:631" *)
  wire _1991_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:634" *)
  wire _1992_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:636" *)
  wire _1993_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:639" *)
  wire _1994_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:641" *)
  wire _1995_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:644" *)
  wire _1996_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:646" *)
  wire _1997_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:649" *)
  wire _1998_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:651" *)
  wire _1999_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:654" *)
  wire _2000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:656" *)
  wire _2001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:659" *)
  wire _2002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:661" *)
  wire _2003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:664" *)
  wire _2004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:666" *)
  wire _2005_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:669" *)
  wire _2006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:671" *)
  wire _2007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:674" *)
  wire _2008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:676" *)
  wire _2009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:679" *)
  wire _2010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:681" *)
  wire _2011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:684" *)
  wire _2012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:686" *)
  wire _2013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:689" *)
  wire _2014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:691" *)
  wire _2015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:694" *)
  wire _2016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:696" *)
  wire _2017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:699" *)
  wire _2018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:701" *)
  wire _2019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:704" *)
  wire _2020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:706" *)
  wire _2021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:709" *)
  wire _2022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:711" *)
  wire _2023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:714" *)
  wire _2024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:716" *)
  wire _2025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:719" *)
  wire _2026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:721" *)
  wire _2027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:724" *)
  wire _2028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:726" *)
  wire _2029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:729" *)
  wire _2030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:731" *)
  wire _2031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:734" *)
  wire _2032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:736" *)
  wire _2033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:739" *)
  wire _2034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:741" *)
  wire _2035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:744" *)
  wire _2036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:746" *)
  wire _2037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:749" *)
  wire _2038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:751" *)
  wire _2039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:754" *)
  wire _2040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:756" *)
  wire _2041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:759" *)
  wire _2042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:761" *)
  wire _2043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:764" *)
  wire _2044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:766" *)
  wire _2045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:769" *)
  wire _2046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:771" *)
  wire _2047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:774" *)
  wire _2048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:776" *)
  wire _2049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:779" *)
  wire _2050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:781" *)
  wire _2051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:784" *)
  wire _2052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:786" *)
  wire _2053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:789" *)
  wire _2054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:791" *)
  wire _2055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:794" *)
  wire _2056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:796" *)
  wire _2057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:799" *)
  wire _2058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:801" *)
  wire _2059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:804" *)
  wire _2060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:806" *)
  wire _2061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:809" *)
  wire _2062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:811" *)
  wire _2063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:814" *)
  wire _2064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:816" *)
  wire _2065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:819" *)
  wire _2066_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:821" *)
  wire _2067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:824" *)
  wire _2068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:826" *)
  wire _2069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:829" *)
  wire _2070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:831" *)
  wire _2071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:834" *)
  wire _2072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:836" *)
  wire _2073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:839" *)
  wire _2074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:841" *)
  wire _2075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:844" *)
  wire _2076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:846" *)
  wire _2077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:849" *)
  wire _2078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:851" *)
  wire _2079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:854" *)
  wire _2080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:856" *)
  wire _2081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:859" *)
  wire _2082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:861" *)
  wire _2083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:864" *)
  wire _2084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:866" *)
  wire _2085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:869" *)
  wire _2086_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:871" *)
  wire _2087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:874" *)
  wire _2088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:876" *)
  wire _2089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:879" *)
  wire _2090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:881" *)
  wire _2091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:884" *)
  wire _2092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:886" *)
  wire _2093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:889" *)
  wire _2094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:891" *)
  wire _2095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:894" *)
  wire _2096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:896" *)
  wire _2097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:899" *)
  wire _2098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:901" *)
  wire _2099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:904" *)
  wire _2100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:906" *)
  wire _2101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:909" *)
  wire _2102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:911" *)
  wire _2103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:914" *)
  wire _2104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:916" *)
  wire _2105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:919" *)
  wire _2106_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:921" *)
  wire _2107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:924" *)
  wire _2108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:926" *)
  wire _2109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:929" *)
  wire _2110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:931" *)
  wire _2111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:934" *)
  wire _2112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:936" *)
  wire _2113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:939" *)
  wire _2114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:941" *)
  wire _2115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:944" *)
  wire _2116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:946" *)
  wire _2117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:949" *)
  wire _2118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:951" *)
  wire _2119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:954" *)
  wire _2120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:956" *)
  wire _2121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:959" *)
  wire _2122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:961" *)
  wire _2123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:964" *)
  wire _2124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:966" *)
  wire _2125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:969" *)
  wire _2126_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:971" *)
  wire _2127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:974" *)
  wire _2128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:976" *)
  wire _2129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:979" *)
  wire _2130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:981" *)
  wire _2131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:984" *)
  wire _2132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:986" *)
  wire _2133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:989" *)
  wire _2134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:991" *)
  wire _2135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:994" *)
  wire _2136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:996" *)
  wire _2137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:999" *)
  wire _2138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:125" *)
  wire _2139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _2140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _2141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *)
  wire _2142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *)
  wire _2143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _2144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _2145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _2146_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _2147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _2148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _2149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *)
  wire _2150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *)
  wire _2151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _2152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _2153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _2154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _2155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _2156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _2157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *)
  wire _2158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *)
  wire _2159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _2160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _2161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _2162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _2163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _2164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _2165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *)
  wire _2166_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *)
  wire _2167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _2168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _2169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _2170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _2171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _2172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _2173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *)
  wire _2174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *)
  wire _2175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _2176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _2177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _2178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _2179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _2180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _2181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *)
  wire _2182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *)
  wire _2183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _2184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _2185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _2186_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _2187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _2188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _2189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *)
  wire _2190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *)
  wire _2191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _2192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _2193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _2194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _2195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _2196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _2197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *)
  wire _2198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *)
  wire _2199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _2200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _2201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _2202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _2203_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _2204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _2205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *)
  wire _2206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *)
  wire _2207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _2208_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _2209_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _2210_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _2211_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _2212_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _2213_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *)
  wire _2214_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *)
  wire _2215_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _2216_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _2217_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _2218_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _2219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *)
  wire _2220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *)
  wire _2221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *)
  wire _2222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *)
  wire _2223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *)
  wire _2224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *)
  wire _2225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *)
  wire _2226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *)
  wire _2227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *)
  wire _2228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *)
  wire _2229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *)
  wire _2230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:211" *)
  wire _2231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2264" *)
  wire _2232_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *)
  wire _2233_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *)
  wire _2234_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *)
  wire _2235_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *)
  wire _2236_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *)
  wire _2237_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *)
  wire _2238_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *)
  wire _2239_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *)
  wire _2240_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *)
  wire _2241_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *)
  wire _2242_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _2243_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *)
  wire _2244_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *)
  wire _2245_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *)
  wire _2246_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *)
  wire _2247_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *)
  wire _2248_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *)
  wire _2249_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *)
  wire _2250_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *)
  wire _2251_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *)
  wire _2252_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _2253_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _2254_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _2255_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *)
  wire _2256_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *)
  wire _2257_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _2258_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *)
  wire _2259_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _2260_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *)
  wire _2261_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *)
  wire _2262_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *)
  wire _2263_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *)
  wire _2264_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *)
  wire _2265_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *)
  wire _2266_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *)
  wire _2267_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *)
  wire _2268_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *)
  wire _2269_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _2270_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _2271_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _2272_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *)
  wire _2273_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *)
  wire _2274_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _2275_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *)
  wire _2276_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _2277_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *)
  wire _2278_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *)
  wire _2279_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *)
  wire _2280_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *)
  wire _2281_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *)
  wire _2282_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *)
  wire _2283_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *)
  wire _2284_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *)
  wire _2285_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *)
  wire _2286_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _2287_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _2288_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _2289_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *)
  wire _2290_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *)
  wire _2291_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _2292_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *)
  wire _2293_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _2294_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *)
  wire _2295_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *)
  wire _2296_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *)
  wire _2297_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *)
  wire _2298_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *)
  wire _2299_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *)
  wire _2300_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *)
  wire _2301_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *)
  wire _2302_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *)
  wire _2303_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _2304_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _2305_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _2306_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *)
  wire _2307_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *)
  wire _2308_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _2309_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *)
  wire _2310_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _2311_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *)
  wire _2312_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *)
  wire _2313_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *)
  wire _2314_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *)
  wire _2315_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *)
  wire _2316_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *)
  wire _2317_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *)
  wire _2318_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *)
  wire _2319_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *)
  wire _2320_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _2321_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _2322_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _2323_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *)
  wire _2324_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *)
  wire _2325_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _2326_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *)
  wire _2327_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _2328_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *)
  wire _2329_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *)
  wire _2330_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *)
  wire _2331_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *)
  wire _2332_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *)
  wire _2333_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *)
  wire _2334_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *)
  wire _2335_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *)
  wire _2336_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *)
  wire _2337_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _2338_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _2339_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _2340_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *)
  wire _2341_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *)
  wire _2342_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _2343_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *)
  wire _2344_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _2345_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *)
  wire _2346_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *)
  wire _2347_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *)
  wire _2348_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *)
  wire _2349_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *)
  wire _2350_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *)
  wire _2351_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *)
  wire _2352_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *)
  wire _2353_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *)
  wire _2354_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _2355_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _2356_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _2357_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *)
  wire _2358_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *)
  wire _2359_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _2360_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *)
  wire _2361_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _2362_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *)
  wire _2363_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *)
  wire _2364_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *)
  wire _2365_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *)
  wire _2366_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *)
  wire _2367_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *)
  wire _2368_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *)
  wire _2369_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *)
  wire _2370_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *)
  wire _2371_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _2372_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _2373_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _2374_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *)
  wire _2375_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *)
  wire _2376_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _2377_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *)
  wire _2378_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _2379_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *)
  wire _2380_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *)
  wire _2381_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *)
  wire _2382_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *)
  wire _2383_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *)
  wire _2384_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *)
  wire _2385_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *)
  wire _2386_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *)
  wire _2387_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *)
  wire _2388_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _2389_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _2390_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _2391_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *)
  wire _2392_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *)
  wire _2393_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _2394_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *)
  wire _2395_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _2396_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *)
  wire _2397_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *)
  wire _2398_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *)
  wire _2399_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *)
  wire _2400_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *)
  wire _2401_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *)
  wire _2402_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *)
  wire _2403_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *)
  wire _2404_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *)
  wire _2405_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _2406_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _2407_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _2408_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *)
  wire _2409_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *)
  wire _2410_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _2411_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *)
  wire _2412_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2413_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2414_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2415_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2416_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2417_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2418_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2419_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *)
  wire _2420_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2421_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2422_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2423_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2424_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2425_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2426_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2427_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2428_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2429_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2430_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2431_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2432_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2433_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2434_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2435_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2436_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2437_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2438_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2439_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2440_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2441_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2442_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2443_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2444_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2445_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *)
  wire _2446_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2457" *)
  wire _2447_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2458" *)
  wire _2448_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2459" *)
  wire _2449_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2460" *)
  wire _2450_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2461" *)
  wire _2451_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2462" *)
  wire _2452_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2463" *)
  wire _2453_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2464" *)
  wire _2454_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2465" *)
  wire _2455_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2466" *)
  wire _2456_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *)
  wire _2457_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *)
  wire _2458_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *)
  wire _2459_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *)
  wire _2460_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *)
  wire _2461_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *)
  wire _2462_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *)
  wire _2463_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *)
  wire _2464_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *)
  wire _2465_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *)
  wire _2466_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *)
  wire _2467_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *)
  wire _2468_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *)
  wire _2469_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *)
  wire _2470_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *)
  wire _2471_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *)
  wire _2472_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *)
  wire _2473_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *)
  wire _2474_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *)
  wire _2475_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *)
  wire _2476_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2477_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *)
  wire _2478_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2633" *)
  wire _2479_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2729" *)
  wire _2480_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2825" *)
  wire _2481_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2921" *)
  wire _2482_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3017" *)
  wire _2483_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3113" *)
  wire _2484_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3209" *)
  wire _2485_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3305" *)
  wire _2486_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3401" *)
  wire _2487_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3497" *)
  wire _2488_;
  wire [6:0] _2489_;
  wire [6:0] _2490_;
  wire [6:0] _2491_;
  wire [6:0] _2492_;
  wire [6:0] _2493_;
  wire [6:0] _2494_;
  wire [6:0] _2495_;
  wire [6:0] _2496_;
  wire [6:0] _2497_;
  wire [6:0] _2498_;
  wire [6:0] _2499_;
  wire [6:0] _2500_;
  wire [6:0] _2501_;
  wire [6:0] _2502_;
  wire [6:0] _2503_;
  wire [6:0] _2504_;
  wire [6:0] _2505_;
  wire [6:0] _2506_;
  wire [6:0] _2507_;
  wire [6:0] _2508_;
  wire [7:0] _2509_;
  wire [7:0] _2510_;
  wire [7:0] _2511_;
  wire [7:0] _2512_;
  wire [7:0] _2513_;
  wire [7:0] _2514_;
  wire [7:0] _2515_;
  wire [7:0] _2516_;
  wire [7:0] _2517_;
  wire [7:0] _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:126" *)
  wire [8:0] _2530_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2115" *)
  wire [8:0] _2531_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2118" *)
  wire [8:0] _2532_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2121" *)
  wire [8:0] _2533_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2124" *)
  wire [8:0] _2534_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2127" *)
  wire [8:0] _2535_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2130" *)
  wire [8:0] _2536_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2133" *)
  wire [8:0] _2537_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2136" *)
  wire [8:0] _2538_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2139" *)
  wire [8:0] _2539_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2142" *)
  wire [8:0] _2540_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2114" *)
  wire [8:0] _2541_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2115" *)
  wire [8:0] _2542_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2117" *)
  wire [8:0] _2543_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2118" *)
  wire [8:0] _2544_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2120" *)
  wire [8:0] _2545_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2121" *)
  wire [8:0] _2546_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2123" *)
  wire [8:0] _2547_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2124" *)
  wire [8:0] _2548_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2126" *)
  wire [8:0] _2549_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2127" *)
  wire [8:0] _2550_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2129" *)
  wire [8:0] _2551_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2130" *)
  wire [8:0] _2552_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2132" *)
  wire [8:0] _2553_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2133" *)
  wire [8:0] _2554_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2135" *)
  wire [8:0] _2555_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2136" *)
  wire [8:0] _2556_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2138" *)
  wire [8:0] _2557_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2139" *)
  wire [8:0] _2558_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2141" *)
  wire [8:0] _2559_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2142" *)
  wire [8:0] _2560_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2491" *)
  wire [7:0] _2561_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2492" *)
  wire [7:0] _2562_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2493" *)
  wire [7:0] _2563_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2494" *)
  wire [7:0] _2564_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2495" *)
  wire [7:0] _2565_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2496" *)
  wire [7:0] _2566_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2497" *)
  wire [7:0] _2567_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2498" *)
  wire [7:0] _2568_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2499" *)
  wire [7:0] _2569_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2500" *)
  wire [7:0] _2570_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2570" *)
  wire [6:0] _2571_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2582" *)
  wire [6:0] _2572_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *)
  wire _2573_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2666" *)
  wire [6:0] _2574_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2678" *)
  wire [6:0] _2575_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *)
  wire _2576_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2762" *)
  wire [6:0] _2577_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2774" *)
  wire [6:0] _2578_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *)
  wire _2579_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2858" *)
  wire [6:0] _2580_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2870" *)
  wire [6:0] _2581_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *)
  wire _2582_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2954" *)
  wire [6:0] _2583_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2966" *)
  wire [6:0] _2584_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *)
  wire _2585_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3050" *)
  wire [6:0] _2586_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3062" *)
  wire [6:0] _2587_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *)
  wire _2588_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3146" *)
  wire [6:0] _2589_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3158" *)
  wire [6:0] _2590_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *)
  wire _2591_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3242" *)
  wire [6:0] _2592_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3254" *)
  wire [6:0] _2593_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *)
  wire _2594_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3338" *)
  wire [6:0] _2595_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3350" *)
  wire [6:0] _2596_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *)
  wire _2597_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3434" *)
  wire [6:0] _2598_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3446" *)
  wire [6:0] _2599_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *)
  wire _2600_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2090" *)
  wire [7:0] adr_ram_rd_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2091" *)
  wire [7:0] adr_ram_rd_data;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2092" *)
  wire adr_ram_rd_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2087" *)
  wire [7:0] adr_ram_wr_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2088" *)
  wire [7:0] adr_ram_wr_data;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2089" *)
  wire adr_ram_wr_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2617" *)
  reg [8:0] cq_rd0_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2618" *)
  reg cq_rd0_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2621" *)
  wire [8:0] cq_rd0_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2619" *)
  wire [8:0] cq_rd0_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2620" *)
  wire [8:0] cq_rd0_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:66" *)
  output [6:0] cq_rd0_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:64" *)
  input cq_rd0_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2558" *)
  reg cq_rd0_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:65" *)
  output cq_rd0_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2713" *)
  reg [8:0] cq_rd1_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2714" *)
  reg cq_rd1_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2717" *)
  wire [8:0] cq_rd1_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2715" *)
  wire [8:0] cq_rd1_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2716" *)
  wire [8:0] cq_rd1_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:69" *)
  output [6:0] cq_rd1_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:67" *)
  input cq_rd1_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2654" *)
  reg cq_rd1_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:68" *)
  output cq_rd1_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2809" *)
  reg [8:0] cq_rd2_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2810" *)
  reg cq_rd2_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2813" *)
  wire [8:0] cq_rd2_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2811" *)
  wire [8:0] cq_rd2_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2812" *)
  wire [8:0] cq_rd2_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:72" *)
  output [6:0] cq_rd2_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:70" *)
  input cq_rd2_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2750" *)
  reg cq_rd2_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:71" *)
  output cq_rd2_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2905" *)
  reg [8:0] cq_rd3_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2906" *)
  reg cq_rd3_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2909" *)
  wire [8:0] cq_rd3_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2907" *)
  wire [8:0] cq_rd3_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2908" *)
  wire [8:0] cq_rd3_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:75" *)
  output [6:0] cq_rd3_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:73" *)
  input cq_rd3_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2846" *)
  reg cq_rd3_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:74" *)
  output cq_rd3_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3001" *)
  reg [8:0] cq_rd4_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3002" *)
  reg cq_rd4_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3005" *)
  wire [8:0] cq_rd4_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3003" *)
  wire [8:0] cq_rd4_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3004" *)
  wire [8:0] cq_rd4_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:78" *)
  output [6:0] cq_rd4_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:76" *)
  input cq_rd4_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2942" *)
  reg cq_rd4_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:77" *)
  output cq_rd4_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3097" *)
  reg [8:0] cq_rd5_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3098" *)
  reg cq_rd5_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3101" *)
  wire [8:0] cq_rd5_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3099" *)
  wire [8:0] cq_rd5_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3100" *)
  wire [8:0] cq_rd5_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:81" *)
  output [6:0] cq_rd5_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:79" *)
  input cq_rd5_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3038" *)
  reg cq_rd5_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:80" *)
  output cq_rd5_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3193" *)
  reg [8:0] cq_rd6_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3194" *)
  reg cq_rd6_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3197" *)
  wire [8:0] cq_rd6_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3195" *)
  wire [8:0] cq_rd6_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3196" *)
  wire [8:0] cq_rd6_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:84" *)
  output [6:0] cq_rd6_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:82" *)
  input cq_rd6_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3134" *)
  reg cq_rd6_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:83" *)
  output cq_rd6_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3289" *)
  reg [8:0] cq_rd7_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3290" *)
  reg cq_rd7_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3293" *)
  wire [8:0] cq_rd7_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3291" *)
  wire [8:0] cq_rd7_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3292" *)
  wire [8:0] cq_rd7_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:87" *)
  output [6:0] cq_rd7_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:85" *)
  input cq_rd7_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3230" *)
  reg cq_rd7_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:86" *)
  output cq_rd7_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3385" *)
  reg [8:0] cq_rd8_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3386" *)
  reg cq_rd8_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3389" *)
  wire [8:0] cq_rd8_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3387" *)
  wire [8:0] cq_rd8_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3388" *)
  wire [8:0] cq_rd8_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:90" *)
  output [6:0] cq_rd8_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:88" *)
  input cq_rd8_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3326" *)
  reg cq_rd8_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:89" *)
  output cq_rd8_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3481" *)
  reg [8:0] cq_rd9_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3482" *)
  reg cq_rd9_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3485" *)
  wire [8:0] cq_rd9_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3483" *)
  wire [8:0] cq_rd9_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3484" *)
  wire [8:0] cq_rd9_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:93" *)
  output [6:0] cq_rd9_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:91" *)
  input cq_rd9_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3422" *)
  reg cq_rd9_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:92" *)
  output cq_rd9_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:180" *)
  wire [7:0] cq_rd_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:181" *)
  wire [7:0] cq_rd_adr_p;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2093" *)
  reg [8:0] cq_rd_count0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2095" *)
  reg [8:0] cq_rd_count1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2097" *)
  reg [8:0] cq_rd_count2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2099" *)
  reg [8:0] cq_rd_count3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2101" *)
  reg [8:0] cq_rd_count4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2103" *)
  reg [8:0] cq_rd_count5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2105" *)
  reg [8:0] cq_rd_count6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2107" *)
  reg [8:0] cq_rd_count7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2109" *)
  reg [8:0] cq_rd_count8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2111" *)
  reg [8:0] cq_rd_count9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2005" *)
  reg [9:0] cq_rd_credit;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:98" *)
  wire [6:0] cq_rd_pd_p;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:97" *)
  wire cq_rd_take;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2549" *)
  wire [9:0] cq_rd_take_elig;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:99" *)
  wire [3:0] cq_rd_take_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3512" *)
  wire [9:0] cq_rd_take_thread_id_is_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3523" *)
  wire [9:0] cq_rd_take_thread_id_is_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3534" *)
  wire [9:0] cq_rd_take_thread_id_is_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3545" *)
  wire [9:0] cq_rd_take_thread_id_is_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3556" *)
  wire [9:0] cq_rd_take_thread_id_is_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3567" *)
  wire [9:0] cq_rd_take_thread_id_is_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3578" *)
  wire [9:0] cq_rd_take_thread_id_is_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3589" *)
  wire [9:0] cq_rd_take_thread_id_is_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3600" *)
  wire [9:0] cq_rd_take_thread_id_is_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3511" *)
  reg [3:0] cq_rd_take_thread_id_last;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:179" *)
  wire [7:0] cq_wr_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:120" *)
  reg cq_wr_busy_int;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:143" *)
  wire cq_wr_busy_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:124" *)
  reg [8:0] cq_wr_count;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:63" *)
  input [6:0] cq_wr_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:57" *)
  output cq_wr_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:58" *)
  input cq_wr_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:59" *)
  input [3:0] cq_wr_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1500" *)
  wire flag_l0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1501" *)
  wire flag_l0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1510" *)
  wire flag_l0_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1600" *)
  wire flag_l0_100;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1601" *)
  wire flag_l0_101;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1602" *)
  wire flag_l0_102;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1603" *)
  wire flag_l0_103;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1604" *)
  wire flag_l0_104;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1605" *)
  wire flag_l0_105;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1606" *)
  wire flag_l0_106;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1607" *)
  wire flag_l0_107;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1608" *)
  wire flag_l0_108;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1609" *)
  wire flag_l0_109;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1511" *)
  wire flag_l0_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1610" *)
  wire flag_l0_110;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1611" *)
  wire flag_l0_111;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1612" *)
  wire flag_l0_112;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1613" *)
  wire flag_l0_113;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1614" *)
  wire flag_l0_114;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1615" *)
  wire flag_l0_115;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1616" *)
  wire flag_l0_116;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1617" *)
  wire flag_l0_117;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1618" *)
  wire flag_l0_118;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1619" *)
  wire flag_l0_119;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1512" *)
  wire flag_l0_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1620" *)
  wire flag_l0_120;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1621" *)
  wire flag_l0_121;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1622" *)
  wire flag_l0_122;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1623" *)
  wire flag_l0_123;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1624" *)
  wire flag_l0_124;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1625" *)
  wire flag_l0_125;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1626" *)
  wire flag_l0_126;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1513" *)
  wire flag_l0_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1514" *)
  wire flag_l0_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1515" *)
  wire flag_l0_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1516" *)
  wire flag_l0_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1517" *)
  wire flag_l0_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1518" *)
  wire flag_l0_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1519" *)
  wire flag_l0_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1502" *)
  wire flag_l0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1520" *)
  wire flag_l0_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1521" *)
  wire flag_l0_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1522" *)
  wire flag_l0_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1523" *)
  wire flag_l0_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1524" *)
  wire flag_l0_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1525" *)
  wire flag_l0_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1526" *)
  wire flag_l0_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1527" *)
  wire flag_l0_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1528" *)
  wire flag_l0_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1529" *)
  wire flag_l0_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1503" *)
  wire flag_l0_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1530" *)
  wire flag_l0_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1531" *)
  wire flag_l0_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1532" *)
  wire flag_l0_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1533" *)
  wire flag_l0_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1534" *)
  wire flag_l0_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1535" *)
  wire flag_l0_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1536" *)
  wire flag_l0_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1537" *)
  wire flag_l0_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1538" *)
  wire flag_l0_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1539" *)
  wire flag_l0_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1504" *)
  wire flag_l0_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1540" *)
  wire flag_l0_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1541" *)
  wire flag_l0_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1542" *)
  wire flag_l0_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1543" *)
  wire flag_l0_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1544" *)
  wire flag_l0_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1545" *)
  wire flag_l0_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1546" *)
  wire flag_l0_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1547" *)
  wire flag_l0_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1548" *)
  wire flag_l0_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1549" *)
  wire flag_l0_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1505" *)
  wire flag_l0_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1550" *)
  wire flag_l0_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1551" *)
  wire flag_l0_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1552" *)
  wire flag_l0_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1553" *)
  wire flag_l0_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1554" *)
  wire flag_l0_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1555" *)
  wire flag_l0_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1556" *)
  wire flag_l0_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1557" *)
  wire flag_l0_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1558" *)
  wire flag_l0_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1559" *)
  wire flag_l0_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1506" *)
  wire flag_l0_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1560" *)
  wire flag_l0_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1561" *)
  wire flag_l0_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1562" *)
  wire flag_l0_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1563" *)
  wire flag_l0_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1564" *)
  wire flag_l0_64;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1565" *)
  wire flag_l0_65;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1566" *)
  wire flag_l0_66;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1567" *)
  wire flag_l0_67;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1568" *)
  wire flag_l0_68;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1569" *)
  wire flag_l0_69;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1507" *)
  wire flag_l0_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1570" *)
  wire flag_l0_70;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1571" *)
  wire flag_l0_71;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1572" *)
  wire flag_l0_72;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1573" *)
  wire flag_l0_73;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1574" *)
  wire flag_l0_74;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1575" *)
  wire flag_l0_75;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1576" *)
  wire flag_l0_76;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1577" *)
  wire flag_l0_77;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1578" *)
  wire flag_l0_78;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1579" *)
  wire flag_l0_79;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1508" *)
  wire flag_l0_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1580" *)
  wire flag_l0_80;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1581" *)
  wire flag_l0_81;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1582" *)
  wire flag_l0_82;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1583" *)
  wire flag_l0_83;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1584" *)
  wire flag_l0_84;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1585" *)
  wire flag_l0_85;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1586" *)
  wire flag_l0_86;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1587" *)
  wire flag_l0_87;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1588" *)
  wire flag_l0_88;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1589" *)
  wire flag_l0_89;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1509" *)
  wire flag_l0_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1590" *)
  wire flag_l0_90;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1591" *)
  wire flag_l0_91;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1592" *)
  wire flag_l0_92;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1593" *)
  wire flag_l0_93;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1594" *)
  wire flag_l0_94;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1595" *)
  wire flag_l0_95;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1596" *)
  wire flag_l0_96;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1597" *)
  wire flag_l0_97;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1598" *)
  wire flag_l0_98;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1599" *)
  wire flag_l0_99;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1627" *)
  wire flag_l1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1628" *)
  wire flag_l1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1637" *)
  wire flag_l1_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1638" *)
  wire flag_l1_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1639" *)
  wire flag_l1_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1640" *)
  wire flag_l1_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1641" *)
  wire flag_l1_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1642" *)
  wire flag_l1_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1643" *)
  wire flag_l1_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1644" *)
  wire flag_l1_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1645" *)
  wire flag_l1_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1646" *)
  wire flag_l1_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1629" *)
  wire flag_l1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1647" *)
  wire flag_l1_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1648" *)
  wire flag_l1_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1649" *)
  wire flag_l1_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1650" *)
  wire flag_l1_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1651" *)
  wire flag_l1_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1652" *)
  wire flag_l1_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1653" *)
  wire flag_l1_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1654" *)
  wire flag_l1_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1655" *)
  wire flag_l1_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1656" *)
  wire flag_l1_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1630" *)
  wire flag_l1_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1657" *)
  wire flag_l1_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1658" *)
  wire flag_l1_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1659" *)
  wire flag_l1_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1660" *)
  wire flag_l1_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1661" *)
  wire flag_l1_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1662" *)
  wire flag_l1_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1663" *)
  wire flag_l1_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1664" *)
  wire flag_l1_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1665" *)
  wire flag_l1_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1666" *)
  wire flag_l1_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1631" *)
  wire flag_l1_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1667" *)
  wire flag_l1_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1668" *)
  wire flag_l1_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1669" *)
  wire flag_l1_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1670" *)
  wire flag_l1_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1671" *)
  wire flag_l1_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1672" *)
  wire flag_l1_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1673" *)
  wire flag_l1_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1674" *)
  wire flag_l1_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1675" *)
  wire flag_l1_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1676" *)
  wire flag_l1_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1632" *)
  wire flag_l1_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1677" *)
  wire flag_l1_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1678" *)
  wire flag_l1_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1679" *)
  wire flag_l1_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1680" *)
  wire flag_l1_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1681" *)
  wire flag_l1_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1682" *)
  wire flag_l1_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1683" *)
  wire flag_l1_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1684" *)
  wire flag_l1_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1685" *)
  wire flag_l1_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1686" *)
  wire flag_l1_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1633" *)
  wire flag_l1_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1687" *)
  wire flag_l1_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1688" *)
  wire flag_l1_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1689" *)
  wire flag_l1_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1634" *)
  wire flag_l1_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1635" *)
  wire flag_l1_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1636" *)
  wire flag_l1_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1690" *)
  wire flag_l2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1691" *)
  wire flag_l2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1700" *)
  wire flag_l2_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1701" *)
  wire flag_l2_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1702" *)
  wire flag_l2_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1703" *)
  wire flag_l2_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1704" *)
  wire flag_l2_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1705" *)
  wire flag_l2_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1706" *)
  wire flag_l2_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1707" *)
  wire flag_l2_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1708" *)
  wire flag_l2_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1709" *)
  wire flag_l2_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1692" *)
  wire flag_l2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1710" *)
  wire flag_l2_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1711" *)
  wire flag_l2_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1712" *)
  wire flag_l2_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1713" *)
  wire flag_l2_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1714" *)
  wire flag_l2_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1715" *)
  wire flag_l2_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1716" *)
  wire flag_l2_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1717" *)
  wire flag_l2_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1718" *)
  wire flag_l2_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1719" *)
  wire flag_l2_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1693" *)
  wire flag_l2_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1720" *)
  wire flag_l2_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1694" *)
  wire flag_l2_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1695" *)
  wire flag_l2_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1696" *)
  wire flag_l2_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1697" *)
  wire flag_l2_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1698" *)
  wire flag_l2_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1699" *)
  wire flag_l2_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1721" *)
  wire flag_l3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1722" *)
  wire flag_l3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1731" *)
  wire flag_l3_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1732" *)
  wire flag_l3_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1733" *)
  wire flag_l3_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1734" *)
  wire flag_l3_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1735" *)
  wire flag_l3_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1723" *)
  wire flag_l3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1724" *)
  wire flag_l3_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1725" *)
  wire flag_l3_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1726" *)
  wire flag_l3_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1727" *)
  wire flag_l3_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1728" *)
  wire flag_l3_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1729" *)
  wire flag_l3_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1730" *)
  wire flag_l3_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1736" *)
  wire flag_l4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1737" *)
  wire flag_l4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1738" *)
  wire flag_l4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1739" *)
  wire flag_l4_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1740" *)
  wire flag_l4_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1741" *)
  wire flag_l4_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1742" *)
  wire flag_l4_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1743" *)
  wire flag_l5_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1744" *)
  wire flag_l5_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1745" *)
  wire flag_l5_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1746" *)
  wire flag_l6_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:203" *)
  wire [7:0] free_adr_index;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:205" *)
  reg [254:0] free_adr_mask;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:204" *)
  wire [254:0] free_adr_mask_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2047" *)
  reg [7:0] head0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2049" *)
  reg [7:0] head1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2051" *)
  reg [7:0] head2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2053" *)
  reg [7:0] head3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2055" *)
  reg [7:0] head4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2057" *)
  reg [7:0] head5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2059" *)
  reg [7:0] head6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2061" *)
  reg [7:0] head7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2063" *)
  reg [7:0] head8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2065" *)
  reg [7:0] head9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1747" *)
  wire index_l0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1748" *)
  wire index_l0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1757" *)
  wire index_l0_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1847" *)
  wire index_l0_100;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1848" *)
  wire index_l0_101;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1849" *)
  wire index_l0_102;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1850" *)
  wire index_l0_103;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1851" *)
  wire index_l0_104;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1852" *)
  wire index_l0_105;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1853" *)
  wire index_l0_106;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1854" *)
  wire index_l0_107;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1855" *)
  wire index_l0_108;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1856" *)
  wire index_l0_109;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1758" *)
  wire index_l0_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1857" *)
  wire index_l0_110;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1858" *)
  wire index_l0_111;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1859" *)
  wire index_l0_112;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1860" *)
  wire index_l0_113;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1861" *)
  wire index_l0_114;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1862" *)
  wire index_l0_115;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1863" *)
  wire index_l0_116;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1864" *)
  wire index_l0_117;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1865" *)
  wire index_l0_118;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1866" *)
  wire index_l0_119;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1759" *)
  wire index_l0_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1867" *)
  wire index_l0_120;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1868" *)
  wire index_l0_121;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1869" *)
  wire index_l0_122;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1870" *)
  wire index_l0_123;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1871" *)
  wire index_l0_124;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1872" *)
  wire index_l0_125;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1873" *)
  wire index_l0_126;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1874" *)
  wire index_l0_127;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1760" *)
  wire index_l0_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1761" *)
  wire index_l0_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1762" *)
  wire index_l0_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1763" *)
  wire index_l0_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1764" *)
  wire index_l0_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1765" *)
  wire index_l0_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1766" *)
  wire index_l0_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1749" *)
  wire index_l0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1767" *)
  wire index_l0_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1768" *)
  wire index_l0_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1769" *)
  wire index_l0_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1770" *)
  wire index_l0_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1771" *)
  wire index_l0_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1772" *)
  wire index_l0_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1773" *)
  wire index_l0_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1774" *)
  wire index_l0_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1775" *)
  wire index_l0_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1776" *)
  wire index_l0_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1750" *)
  wire index_l0_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1777" *)
  wire index_l0_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1778" *)
  wire index_l0_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1779" *)
  wire index_l0_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1780" *)
  wire index_l0_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1781" *)
  wire index_l0_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1782" *)
  wire index_l0_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1783" *)
  wire index_l0_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1784" *)
  wire index_l0_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1785" *)
  wire index_l0_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1786" *)
  wire index_l0_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1751" *)
  wire index_l0_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1787" *)
  wire index_l0_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1788" *)
  wire index_l0_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1789" *)
  wire index_l0_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1790" *)
  wire index_l0_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1791" *)
  wire index_l0_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1792" *)
  wire index_l0_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1793" *)
  wire index_l0_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1794" *)
  wire index_l0_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1795" *)
  wire index_l0_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1796" *)
  wire index_l0_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1752" *)
  wire index_l0_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1797" *)
  wire index_l0_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1798" *)
  wire index_l0_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1799" *)
  wire index_l0_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1800" *)
  wire index_l0_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1801" *)
  wire index_l0_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1802" *)
  wire index_l0_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1803" *)
  wire index_l0_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1804" *)
  wire index_l0_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1805" *)
  wire index_l0_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1806" *)
  wire index_l0_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1753" *)
  wire index_l0_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1807" *)
  wire index_l0_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1808" *)
  wire index_l0_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1809" *)
  wire index_l0_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1810" *)
  wire index_l0_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1811" *)
  wire index_l0_64;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1812" *)
  wire index_l0_65;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1813" *)
  wire index_l0_66;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1814" *)
  wire index_l0_67;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1815" *)
  wire index_l0_68;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1816" *)
  wire index_l0_69;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1754" *)
  wire index_l0_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1817" *)
  wire index_l0_70;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1818" *)
  wire index_l0_71;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1819" *)
  wire index_l0_72;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1820" *)
  wire index_l0_73;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1821" *)
  wire index_l0_74;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1822" *)
  wire index_l0_75;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1823" *)
  wire index_l0_76;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1824" *)
  wire index_l0_77;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1825" *)
  wire index_l0_78;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1826" *)
  wire index_l0_79;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1755" *)
  wire index_l0_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1827" *)
  wire index_l0_80;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1828" *)
  wire index_l0_81;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1829" *)
  wire index_l0_82;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1830" *)
  wire index_l0_83;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1831" *)
  wire index_l0_84;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1832" *)
  wire index_l0_85;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1833" *)
  wire index_l0_86;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1834" *)
  wire index_l0_87;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1835" *)
  wire index_l0_88;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1836" *)
  wire index_l0_89;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1756" *)
  wire index_l0_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1837" *)
  wire index_l0_90;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1838" *)
  wire index_l0_91;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1839" *)
  wire index_l0_92;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1840" *)
  wire index_l0_93;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1841" *)
  wire index_l0_94;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1842" *)
  wire index_l0_95;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1843" *)
  wire index_l0_96;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1844" *)
  wire index_l0_97;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1845" *)
  wire index_l0_98;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1846" *)
  wire index_l0_99;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1875" *)
  wire [1:0] index_l1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1876" *)
  wire [1:0] index_l1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1885" *)
  wire [1:0] index_l1_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1886" *)
  wire [1:0] index_l1_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1887" *)
  wire [1:0] index_l1_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1888" *)
  wire [1:0] index_l1_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1889" *)
  wire [1:0] index_l1_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1890" *)
  wire [1:0] index_l1_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1891" *)
  wire [1:0] index_l1_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1892" *)
  wire [1:0] index_l1_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1893" *)
  wire [1:0] index_l1_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1894" *)
  wire [1:0] index_l1_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1877" *)
  wire [1:0] index_l1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1895" *)
  wire [1:0] index_l1_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1896" *)
  wire [1:0] index_l1_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1897" *)
  wire [1:0] index_l1_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1898" *)
  wire [1:0] index_l1_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1899" *)
  wire [1:0] index_l1_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1900" *)
  wire [1:0] index_l1_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1901" *)
  wire [1:0] index_l1_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1902" *)
  wire [1:0] index_l1_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1903" *)
  wire [1:0] index_l1_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1904" *)
  wire [1:0] index_l1_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1878" *)
  wire [1:0] index_l1_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1905" *)
  wire [1:0] index_l1_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1906" *)
  wire [1:0] index_l1_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1907" *)
  wire [1:0] index_l1_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1908" *)
  wire [1:0] index_l1_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1909" *)
  wire [1:0] index_l1_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1910" *)
  wire [1:0] index_l1_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1911" *)
  wire [1:0] index_l1_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1912" *)
  wire [1:0] index_l1_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1913" *)
  wire [1:0] index_l1_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1914" *)
  wire [1:0] index_l1_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1879" *)
  wire [1:0] index_l1_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1915" *)
  wire [1:0] index_l1_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1916" *)
  wire [1:0] index_l1_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1917" *)
  wire [1:0] index_l1_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1918" *)
  wire [1:0] index_l1_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1919" *)
  wire [1:0] index_l1_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1920" *)
  wire [1:0] index_l1_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1921" *)
  wire [1:0] index_l1_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1922" *)
  wire [1:0] index_l1_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1923" *)
  wire [1:0] index_l1_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1924" *)
  wire [1:0] index_l1_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1880" *)
  wire [1:0] index_l1_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1925" *)
  wire [1:0] index_l1_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1926" *)
  wire [1:0] index_l1_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1927" *)
  wire [1:0] index_l1_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1928" *)
  wire [1:0] index_l1_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1929" *)
  wire [1:0] index_l1_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1930" *)
  wire [1:0] index_l1_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1931" *)
  wire [1:0] index_l1_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1932" *)
  wire [1:0] index_l1_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1933" *)
  wire [1:0] index_l1_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1934" *)
  wire [1:0] index_l1_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1881" *)
  wire [1:0] index_l1_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1935" *)
  wire [1:0] index_l1_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1936" *)
  wire [1:0] index_l1_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1937" *)
  wire [1:0] index_l1_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1938" *)
  wire [1:0] index_l1_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1882" *)
  wire [1:0] index_l1_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1883" *)
  wire [1:0] index_l1_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1884" *)
  wire [1:0] index_l1_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1939" *)
  wire [2:0] index_l2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1940" *)
  wire [2:0] index_l2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1949" *)
  wire [2:0] index_l2_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1950" *)
  wire [2:0] index_l2_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1951" *)
  wire [2:0] index_l2_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1952" *)
  wire [2:0] index_l2_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1953" *)
  wire [2:0] index_l2_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1954" *)
  wire [2:0] index_l2_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1955" *)
  wire [2:0] index_l2_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1956" *)
  wire [2:0] index_l2_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1957" *)
  wire [2:0] index_l2_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1958" *)
  wire [2:0] index_l2_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1941" *)
  wire [2:0] index_l2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1959" *)
  wire [2:0] index_l2_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1960" *)
  wire [2:0] index_l2_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1961" *)
  wire [2:0] index_l2_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1962" *)
  wire [2:0] index_l2_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1963" *)
  wire [2:0] index_l2_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1964" *)
  wire [2:0] index_l2_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1965" *)
  wire [2:0] index_l2_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1966" *)
  wire [2:0] index_l2_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1967" *)
  wire [2:0] index_l2_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1968" *)
  wire [2:0] index_l2_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1942" *)
  wire [2:0] index_l2_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1969" *)
  wire [2:0] index_l2_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1970" *)
  wire [2:0] index_l2_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1943" *)
  wire [2:0] index_l2_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1944" *)
  wire [2:0] index_l2_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1945" *)
  wire [2:0] index_l2_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1946" *)
  wire [2:0] index_l2_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1947" *)
  wire [2:0] index_l2_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1948" *)
  wire [2:0] index_l2_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1971" *)
  wire [3:0] index_l3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1972" *)
  wire [3:0] index_l3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1981" *)
  wire [3:0] index_l3_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1982" *)
  wire [3:0] index_l3_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1983" *)
  wire [3:0] index_l3_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1984" *)
  wire [3:0] index_l3_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1985" *)
  wire [3:0] index_l3_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1986" *)
  wire [3:0] index_l3_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1973" *)
  wire [3:0] index_l3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1974" *)
  wire [3:0] index_l3_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1975" *)
  wire [3:0] index_l3_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1976" *)
  wire [3:0] index_l3_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1977" *)
  wire [3:0] index_l3_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1978" *)
  wire [3:0] index_l3_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1979" *)
  wire [3:0] index_l3_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1980" *)
  wire [3:0] index_l3_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1987" *)
  wire [4:0] index_l4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1988" *)
  wire [4:0] index_l4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1989" *)
  wire [4:0] index_l4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1990" *)
  wire [4:0] index_l4_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1991" *)
  wire [4:0] index_l4_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1992" *)
  wire [4:0] index_l4_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1993" *)
  wire [4:0] index_l4_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1994" *)
  wire [4:0] index_l4_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1995" *)
  wire [5:0] index_l5_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1996" *)
  wire [5:0] index_l5_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1997" *)
  wire [5:0] index_l5_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1998" *)
  wire [5:0] index_l5_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1999" *)
  wire [6:0] index_l6_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2000" *)
  wire [6:0] index_l6_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2001" *)
  wire [7:0] index_l7_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:55" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:107" *)
  wire nvdla_core_clk_mgated;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:106" *)
  wire nvdla_core_clk_mgated_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:103" *)
  wire nvdla_core_clk_mgated_skid;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:104" *)
  wire nvdla_core_clk_mgated_skid_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:56" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:94" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2527" *)
  reg [7:0] rd_adr_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2551" *)
  wire rd_bypassing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2647" *)
  wire rd_bypassing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2743" *)
  wire rd_bypassing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2839" *)
  wire rd_bypassing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2935" *)
  wire rd_bypassing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3031" *)
  wire rd_bypassing5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3127" *)
  wire rd_bypassing6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3223" *)
  wire rd_bypassing7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3319" *)
  wire rd_bypassing8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3415" *)
  wire rd_bypassing9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2094" *)
  wire [8:0] rd_count0_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2096" *)
  wire [8:0] rd_count1_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2098" *)
  wire [8:0] rd_count2_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2100" *)
  wire [8:0] rd_count3_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2102" *)
  wire [8:0] rd_count4_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2104" *)
  wire [8:0] rd_count5_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2106" *)
  wire [8:0] rd_count6_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2108" *)
  wire [8:0] rd_count7_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2110" *)
  wire [8:0] rd_count8_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2112" *)
  wire [8:0] rd_count9_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:182" *)
  wire rd_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:194" *)
  wire rd_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:202" *)
  wire [7:0] rd_popping_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2550" *)
  wire rd_pre_bypassing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2646" *)
  wire rd_pre_bypassing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2742" *)
  wire rd_pre_bypassing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2838" *)
  wire rd_pre_bypassing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2934" *)
  wire rd_pre_bypassing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3030" *)
  wire rd_pre_bypassing5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3126" *)
  wire rd_pre_bypassing6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3222" *)
  wire rd_pre_bypassing7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3318" *)
  wire rd_pre_bypassing8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3414" *)
  wire rd_pre_bypassing9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:197" *)
  wire rd_pushing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2027" *)
  wire rd_pushing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2028" *)
  wire rd_pushing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2029" *)
  wire rd_pushing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2030" *)
  wire rd_pushing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2031" *)
  wire rd_pushing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2032" *)
  wire rd_pushing5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2033" *)
  wire rd_pushing6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2034" *)
  wire rd_pushing7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2035" *)
  wire rd_pushing8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2036" *)
  wire rd_pushing9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:199" *)
  wire [7:0] rd_pushing_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2006" *)
  reg rd_pushing_q;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:198" *)
  wire [3:0] rd_pushing_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2552" *)
  reg [6:0] rd_skid0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2555" *)
  reg rd_skid0_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2553" *)
  reg [6:0] rd_skid0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2556" *)
  reg rd_skid0_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2554" *)
  reg [6:0] rd_skid0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2557" *)
  reg rd_skid0_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2648" *)
  reg [6:0] rd_skid1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2651" *)
  reg rd_skid1_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2649" *)
  reg [6:0] rd_skid1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2652" *)
  reg rd_skid1_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2650" *)
  reg [6:0] rd_skid1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2653" *)
  reg rd_skid1_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2744" *)
  reg [6:0] rd_skid2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2747" *)
  reg rd_skid2_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2745" *)
  reg [6:0] rd_skid2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2748" *)
  reg rd_skid2_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2746" *)
  reg [6:0] rd_skid2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2749" *)
  reg rd_skid2_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2840" *)
  reg [6:0] rd_skid3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2843" *)
  reg rd_skid3_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2841" *)
  reg [6:0] rd_skid3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2844" *)
  reg rd_skid3_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2842" *)
  reg [6:0] rd_skid3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2845" *)
  reg rd_skid3_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2936" *)
  reg [6:0] rd_skid4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2939" *)
  reg rd_skid4_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2937" *)
  reg [6:0] rd_skid4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2940" *)
  reg rd_skid4_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2938" *)
  reg [6:0] rd_skid4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2941" *)
  reg rd_skid4_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3032" *)
  reg [6:0] rd_skid5_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3035" *)
  reg rd_skid5_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3033" *)
  reg [6:0] rd_skid5_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3036" *)
  reg rd_skid5_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3034" *)
  reg [6:0] rd_skid5_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3037" *)
  reg rd_skid5_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3128" *)
  reg [6:0] rd_skid6_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3131" *)
  reg rd_skid6_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3129" *)
  reg [6:0] rd_skid6_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3132" *)
  reg rd_skid6_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3130" *)
  reg [6:0] rd_skid6_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3133" *)
  reg rd_skid6_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3224" *)
  reg [6:0] rd_skid7_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3227" *)
  reg rd_skid7_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3225" *)
  reg [6:0] rd_skid7_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3228" *)
  reg rd_skid7_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3226" *)
  reg [6:0] rd_skid7_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3229" *)
  reg rd_skid7_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3320" *)
  reg [6:0] rd_skid8_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3323" *)
  reg rd_skid8_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3321" *)
  reg [6:0] rd_skid8_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3324" *)
  reg rd_skid8_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3322" *)
  reg [6:0] rd_skid8_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3325" *)
  reg rd_skid8_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3416" *)
  reg [6:0] rd_skid9_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3419" *)
  reg rd_skid9_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3417" *)
  reg [6:0] rd_skid9_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3420" *)
  reg rd_skid9_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3418" *)
  reg [6:0] rd_skid9_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3421" *)
  reg rd_skid9_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2037" *)
  wire rd_take0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2038" *)
  wire rd_take1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2039" *)
  wire rd_take2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2040" *)
  wire rd_take3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2041" *)
  wire rd_take4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2042" *)
  wire rd_take5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2043" *)
  wire rd_take6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2044" *)
  wire rd_take7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2045" *)
  wire rd_take8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2046" *)
  wire rd_take9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2525" *)
  reg rd_take_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2068" *)
  wire rd_take_dly_cg;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2067" *)
  reg [9:0] rd_take_n_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2048" *)
  reg [7:0] tail0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2050" *)
  reg [7:0] tail1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2052" *)
  reg [7:0] tail2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2054" *)
  reg [7:0] tail3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2056" *)
  reg [7:0] tail4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2058" *)
  reg [7:0] tail5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2060" *)
  reg [7:0] tail6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2062" *)
  reg [7:0] tail7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2064" *)
  reg [7:0] tail8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2066" *)
  reg [7:0] tail9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2248" *)
  reg [9:0] update_head;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2249" *)
  wire [9:0] update_head_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2069" *)
  wire update_rd_take_n_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:178" *)
  wire wr_adr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:101" *)
  wire wr_bypassing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:128" *)
  wire [8:0] wr_count_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:131" *)
  wire wr_count_next_is_256;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:127" *)
  wire [8:0] wr_count_next_no_wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:130" *)
  wire wr_count_next_no_wr_popping_is_256;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:126" *)
  wire [8:0] wr_count_next_wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:133" *)
  wire [8:0] wr_limit_muxed;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:134" *)
  wire [8:0] wr_limit_reg;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:123" *)
  wire wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:173" *)
  wire wr_pushing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:174" *)
  wire [3:0] wr_pushing_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:119" *)
  wire wr_reserving;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:125" *)
  wire wr_reserving_and_not_bypassing;
  assign _0373_ = cq_wr_count + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:127" *) 1'b1;
  assign _0374_ = cq_rd_count0 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2114" *) 1'b1;
  assign _0375_ = cq_rd_count1 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2117" *) 1'b1;
  assign _0376_ = cq_rd_count2 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2120" *) 1'b1;
  assign _0377_ = cq_rd_count3 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2123" *) 1'b1;
  assign _0378_ = cq_rd_count4 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2126" *) 1'b1;
  assign _0379_ = cq_rd_count5 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2129" *) 1'b1;
  assign _0380_ = cq_rd_count6 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2132" *) 1'b1;
  assign _0381_ = cq_rd_count7 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2135" *) 1'b1;
  assign _0382_ = cq_rd_count8 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2138" *) 1'b1;
  assign _0383_ = cq_rd_count9 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2141" *) 1'b1;
  assign cq_rd0_credits_wo_take_next = cq_rd0_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2619" *) cq_rd_credit[0];
  assign cq_rd1_credits_wo_take_next = cq_rd1_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2715" *) cq_rd_credit[1];
  assign cq_rd2_credits_wo_take_next = cq_rd2_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2811" *) cq_rd_credit[2];
  assign cq_rd3_credits_wo_take_next = cq_rd3_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2907" *) cq_rd_credit[3];
  assign cq_rd4_credits_wo_take_next = cq_rd4_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3003" *) cq_rd_credit[4];
  assign cq_rd5_credits_wo_take_next = cq_rd5_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3099" *) cq_rd_credit[5];
  assign cq_rd6_credits_wo_take_next = cq_rd6_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3195" *) cq_rd_credit[6];
  assign cq_rd7_credits_wo_take_next = cq_rd7_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3291" *) cq_rd_credit[7];
  assign cq_rd8_credits_wo_take_next = cq_rd8_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3387" *) cq_rd_credit[8];
  assign cq_rd9_credits_wo_take_next = cq_rd9_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3483" *) cq_rd_credit[9];
  assign _0384_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1001" *) 8'b10011011;
  assign _0385_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1004" *) 8'b10011100;
  assign _0386_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1006" *) 8'b10011100;
  assign _0387_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1009" *) 8'b10011101;
  assign _0388_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1011" *) 8'b10011101;
  assign _0389_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1014" *) 8'b10011110;
  assign _0390_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1016" *) 8'b10011110;
  assign _0391_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1019" *) 8'b10011111;
  assign _0392_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1021" *) 8'b10011111;
  assign _0393_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1024" *) 8'b10100000;
  assign _0394_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1026" *) 8'b10100000;
  assign _0395_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1029" *) 8'b10100001;
  assign _0396_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1031" *) 8'b10100001;
  assign _0397_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1034" *) 8'b10100010;
  assign _0398_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1036" *) 8'b10100010;
  assign _0399_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1039" *) 8'b10100011;
  assign _0400_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1041" *) 8'b10100011;
  assign _0401_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1044" *) 8'b10100100;
  assign _0402_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1046" *) 8'b10100100;
  assign _0403_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1049" *) 8'b10100101;
  assign _0404_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1051" *) 8'b10100101;
  assign _0405_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1054" *) 8'b10100110;
  assign _0406_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1056" *) 8'b10100110;
  assign _0407_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1059" *) 8'b10100111;
  assign _0408_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1061" *) 8'b10100111;
  assign _0409_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1064" *) 8'b10101000;
  assign _0410_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1066" *) 8'b10101000;
  assign _0411_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1069" *) 8'b10101001;
  assign _0412_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1071" *) 8'b10101001;
  assign _0413_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1074" *) 8'b10101010;
  assign _0414_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1076" *) 8'b10101010;
  assign _0415_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1079" *) 8'b10101011;
  assign _0416_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1081" *) 8'b10101011;
  assign _0417_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1084" *) 8'b10101100;
  assign _0418_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1086" *) 8'b10101100;
  assign _0419_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1089" *) 8'b10101101;
  assign _0420_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1091" *) 8'b10101101;
  assign _0421_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1094" *) 8'b10101110;
  assign _0422_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1096" *) 8'b10101110;
  assign _0423_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1099" *) 8'b10101111;
  assign _0424_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1101" *) 8'b10101111;
  assign _0425_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1104" *) 8'b10110000;
  assign _0426_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1106" *) 8'b10110000;
  assign _0427_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1109" *) 8'b10110001;
  assign _0428_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1111" *) 8'b10110001;
  assign _0429_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1114" *) 8'b10110010;
  assign _0430_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1116" *) 8'b10110010;
  assign _0431_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1119" *) 8'b10110011;
  assign _0432_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1121" *) 8'b10110011;
  assign _0433_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1124" *) 8'b10110100;
  assign _0434_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1126" *) 8'b10110100;
  assign _0435_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1129" *) 8'b10110101;
  assign _0436_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1131" *) 8'b10110101;
  assign _0437_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1134" *) 8'b10110110;
  assign _0438_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1136" *) 8'b10110110;
  assign _0439_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1139" *) 8'b10110111;
  assign _0440_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1141" *) 8'b10110111;
  assign _0441_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1144" *) 8'b10111000;
  assign _0442_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1146" *) 8'b10111000;
  assign _0443_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1149" *) 8'b10111001;
  assign _0444_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1151" *) 8'b10111001;
  assign _0445_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1154" *) 8'b10111010;
  assign _0446_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1156" *) 8'b10111010;
  assign _0447_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1159" *) 8'b10111011;
  assign _0448_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1161" *) 8'b10111011;
  assign _0449_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1164" *) 8'b10111100;
  assign _0450_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1166" *) 8'b10111100;
  assign _0451_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1169" *) 8'b10111101;
  assign _0452_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1171" *) 8'b10111101;
  assign _0453_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1174" *) 8'b10111110;
  assign _0454_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1176" *) 8'b10111110;
  assign _0455_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1179" *) 8'b10111111;
  assign _0456_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1181" *) 8'b10111111;
  assign _0457_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1184" *) 8'b11000000;
  assign _0458_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1186" *) 8'b11000000;
  assign _0459_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1189" *) 8'b11000001;
  assign _0460_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1191" *) 8'b11000001;
  assign _0461_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1194" *) 8'b11000010;
  assign _0462_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1196" *) 8'b11000010;
  assign _0463_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1199" *) 8'b11000011;
  assign _0464_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1201" *) 8'b11000011;
  assign _0465_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1204" *) 8'b11000100;
  assign _0466_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1206" *) 8'b11000100;
  assign _0467_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1209" *) 8'b11000101;
  assign _0468_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1211" *) 8'b11000101;
  assign _0469_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1214" *) 8'b11000110;
  assign _0470_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1216" *) 8'b11000110;
  assign _0471_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1219" *) 8'b11000111;
  assign _0472_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1221" *) 8'b11000111;
  assign _0473_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1224" *) 8'b11001000;
  assign _0474_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1226" *) 8'b11001000;
  assign _0475_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1229" *) 8'b11001001;
  assign _0476_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1231" *) 8'b11001001;
  assign _0477_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1234" *) 8'b11001010;
  assign _0478_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1236" *) 8'b11001010;
  assign _0479_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1239" *) 8'b11001011;
  assign _0480_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1241" *) 8'b11001011;
  assign _0481_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1244" *) 8'b11001100;
  assign _0482_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1246" *) 8'b11001100;
  assign _0483_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1249" *) 8'b11001101;
  assign _0484_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1251" *) 8'b11001101;
  assign _0485_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1254" *) 8'b11001110;
  assign _0486_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1256" *) 8'b11001110;
  assign _0487_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1259" *) 8'b11001111;
  assign _0488_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1261" *) 8'b11001111;
  assign _0489_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1264" *) 8'b11010000;
  assign _0490_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1266" *) 8'b11010000;
  assign _0491_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1269" *) 8'b11010001;
  assign _0492_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1271" *) 8'b11010001;
  assign _0493_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1274" *) 8'b11010010;
  assign _0494_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1276" *) 8'b11010010;
  assign _0495_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1279" *) 8'b11010011;
  assign _0496_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1281" *) 8'b11010011;
  assign _0497_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1284" *) 8'b11010100;
  assign _0498_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1286" *) 8'b11010100;
  assign _0499_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1289" *) 8'b11010101;
  assign _0500_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1291" *) 8'b11010101;
  assign _0501_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1294" *) 8'b11010110;
  assign _0502_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1296" *) 8'b11010110;
  assign _0503_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1299" *) 8'b11010111;
  assign wr_count_next_no_wr_popping_is_256 = wr_count_next_no_wr_popping == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:130" *) 9'b100000000;
  assign _0504_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1301" *) 8'b11010111;
  assign _0505_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1304" *) 8'b11011000;
  assign _0506_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1306" *) 8'b11011000;
  assign _0507_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1309" *) 8'b11011001;
  assign _0508_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1311" *) 8'b11011001;
  assign _0509_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1314" *) 8'b11011010;
  assign _0510_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1316" *) 8'b11011010;
  assign _0511_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1319" *) 8'b11011011;
  assign _0512_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1321" *) 8'b11011011;
  assign _0513_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1324" *) 8'b11011100;
  assign _0514_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1326" *) 8'b11011100;
  assign _0515_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1329" *) 8'b11011101;
  assign _0516_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1331" *) 8'b11011101;
  assign _0517_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1334" *) 8'b11011110;
  assign _0518_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1336" *) 8'b11011110;
  assign _0519_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1339" *) 8'b11011111;
  assign _0520_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1341" *) 8'b11011111;
  assign _0521_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1344" *) 8'b11100000;
  assign _0522_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1346" *) 8'b11100000;
  assign _0523_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1349" *) 8'b11100001;
  assign _0524_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1351" *) 8'b11100001;
  assign _0525_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1354" *) 8'b11100010;
  assign _0526_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1356" *) 8'b11100010;
  assign _0527_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1359" *) 8'b11100011;
  assign _0528_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1361" *) 8'b11100011;
  assign _0529_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1364" *) 8'b11100100;
  assign _0530_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1366" *) 8'b11100100;
  assign _0531_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1369" *) 8'b11100101;
  assign _0532_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1371" *) 8'b11100101;
  assign _0533_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1374" *) 8'b11100110;
  assign _0534_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1376" *) 8'b11100110;
  assign _0535_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1379" *) 8'b11100111;
  assign _0536_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1381" *) 8'b11100111;
  assign _0537_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1384" *) 8'b11101000;
  assign _0538_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1386" *) 8'b11101000;
  assign _0539_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1389" *) 8'b11101001;
  assign _0540_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1391" *) 8'b11101001;
  assign _0541_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1394" *) 8'b11101010;
  assign _0542_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1396" *) 8'b11101010;
  assign _0543_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1399" *) 8'b11101011;
  assign _0544_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1401" *) 8'b11101011;
  assign _0545_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1404" *) 8'b11101100;
  assign _0546_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1406" *) 8'b11101100;
  assign _0547_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1409" *) 8'b11101101;
  assign _0548_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1411" *) 8'b11101101;
  assign _0549_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1414" *) 8'b11101110;
  assign _0550_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1416" *) 8'b11101110;
  assign _0551_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1419" *) 8'b11101111;
  assign _0552_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1421" *) 8'b11101111;
  assign _0553_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1424" *) 8'b11110000;
  assign _0554_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1426" *) 8'b11110000;
  assign _0555_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1429" *) 8'b11110001;
  assign _0556_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1431" *) 8'b11110001;
  assign _0557_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1434" *) 8'b11110010;
  assign _0558_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1436" *) 8'b11110010;
  assign _0559_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1439" *) 8'b11110011;
  assign _0560_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1441" *) 8'b11110011;
  assign _0561_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1444" *) 8'b11110100;
  assign _0562_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1446" *) 8'b11110100;
  assign _0563_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1449" *) 8'b11110101;
  assign _0564_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1451" *) 8'b11110101;
  assign _0565_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1454" *) 8'b11110110;
  assign _0566_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1456" *) 8'b11110110;
  assign _0567_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1459" *) 8'b11110111;
  assign _0568_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1461" *) 8'b11110111;
  assign _0569_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1464" *) 8'b11111000;
  assign _0570_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1466" *) 8'b11111000;
  assign _0571_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1469" *) 8'b11111001;
  assign _0572_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1471" *) 8'b11111001;
  assign _0573_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1474" *) 8'b11111010;
  assign _0574_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1476" *) 8'b11111010;
  assign _0575_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1479" *) 8'b11111011;
  assign _0576_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1481" *) 8'b11111011;
  assign _0577_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1484" *) 8'b11111100;
  assign _0578_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1486" *) 8'b11111100;
  assign _0579_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1489" *) 8'b11111101;
  assign _0580_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1491" *) 8'b11111101;
  assign _0581_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1494" *) 8'b11111110;
  assign _0582_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1496" *) 8'b11111110;
  assign _0583_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2013" *) cq_wr_thread_id;
  assign _0584_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2014" *) 1'b1;
  assign _0585_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2015" *) 2'b10;
  assign _0586_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2016" *) 2'b11;
  assign _0587_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2017" *) 3'b100;
  assign _0588_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2018" *) 3'b101;
  assign _0589_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2019" *) 3'b110;
  assign _0590_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2020" *) 3'b111;
  assign _0591_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2021" *) 4'b1000;
  assign _0592_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2022" *) 4'b1001;
  assign _0593_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2037" *) cq_rd_take_thread_id;
  assign _0594_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2038" *) 1'b1;
  assign _0595_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2039" *) 2'b10;
  assign _0596_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2040" *) 2'b11;
  assign _0597_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2041" *) 3'b100;
  assign _0598_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2042" *) 3'b101;
  assign _0599_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2043" *) 3'b110;
  assign _0600_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2044" *) 3'b111;
  assign _0601_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2045" *) 4'b1000;
  assign _0602_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2046" *) 4'b1001;
  assign _0603_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:224" *) rd_adr_dly;
  assign _0604_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:226" *) adr_ram_wr_data;
  assign _0605_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2285" *) cq_rd_count0;
  assign _0606_ = cq_rd_count0 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *) 1'b1;
  assign _0607_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:229" *) 1'b1;
  assign _0608_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2300" *) cq_rd_count1;
  assign _0609_ = cq_rd_count1 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *) 1'b1;
  assign _0610_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:231" *) 1'b1;
  assign _0611_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2315" *) cq_rd_count2;
  assign _0612_ = cq_rd_count2 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *) 1'b1;
  assign _0613_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2330" *) cq_rd_count3;
  assign _0614_ = cq_rd_count3 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *) 1'b1;
  assign _0615_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:234" *) 2'b10;
  assign _0616_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2345" *) cq_rd_count4;
  assign _0617_ = cq_rd_count4 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *) 1'b1;
  assign _0618_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:236" *) 2'b10;
  assign _0619_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2360" *) cq_rd_count5;
  assign _0620_ = cq_rd_count5 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *) 1'b1;
  assign _0621_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2375" *) cq_rd_count6;
  assign _0622_ = cq_rd_count6 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *) 1'b1;
  assign _0623_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:239" *) 2'b11;
  assign _0624_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2390" *) cq_rd_count7;
  assign _0625_ = cq_rd_count7 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *) 1'b1;
  assign _0626_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2405" *) cq_rd_count8;
  assign _0627_ = cq_rd_count8 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *) 1'b1;
  assign _0628_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:241" *) 2'b11;
  assign _0629_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2420" *) cq_rd_count9;
  assign _0630_ = cq_rd_count9 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *) 1'b1;
  assign _0631_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:244" *) 3'b100;
  assign _0632_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:246" *) 3'b100;
  assign _0633_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:249" *) 3'b101;
  assign _0634_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:251" *) 3'b101;
  assign _0635_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:254" *) 3'b110;
  assign _0636_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:256" *) 3'b110;
  assign _0637_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:259" *) 3'b111;
  assign _0638_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:261" *) 3'b111;
  assign _0639_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) cq_rd0_credits;
  assign _0640_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:264" *) 4'b1000;
  assign _0641_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:266" *) 4'b1000;
  assign _0642_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:269" *) 4'b1001;
  assign _0643_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:271" *) 4'b1001;
  assign _0644_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) cq_rd1_credits;
  assign _0645_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:274" *) 4'b1010;
  assign _0646_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:276" *) 4'b1010;
  assign _0647_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:279" *) 4'b1011;
  assign _0648_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:281" *) 4'b1011;
  assign _0649_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) cq_rd2_credits;
  assign _0650_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:284" *) 4'b1100;
  assign _0651_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:286" *) 4'b1100;
  assign _0652_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:289" *) 4'b1101;
  assign _0653_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:291" *) 4'b1101;
  assign _0654_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) cq_rd3_credits;
  assign _0655_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:294" *) 4'b1110;
  assign _0656_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:296" *) 4'b1110;
  assign _0657_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:299" *) 4'b1111;
  assign _0658_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:301" *) 4'b1111;
  assign _0659_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) cq_rd4_credits;
  assign _0660_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:304" *) 5'b10000;
  assign _0661_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:306" *) 5'b10000;
  assign _0662_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:309" *) 5'b10001;
  assign _0663_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) cq_rd5_credits;
  assign _0664_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:311" *) 5'b10001;
  assign _0665_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:314" *) 5'b10010;
  assign _0666_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:316" *) 5'b10010;
  assign _0667_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:319" *) 5'b10011;
  assign _0668_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) cq_rd6_credits;
  assign _0669_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:321" *) 5'b10011;
  assign _0670_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:324" *) 5'b10100;
  assign _0671_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:326" *) 5'b10100;
  assign _0672_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:329" *) 5'b10101;
  assign _0673_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) cq_rd7_credits;
  assign _0674_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:331" *) 5'b10101;
  assign _0675_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:334" *) 5'b10110;
  assign _0676_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:336" *) 5'b10110;
  assign _0677_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:339" *) 5'b10111;
  assign _0678_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) cq_rd8_credits;
  assign _0679_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:341" *) 5'b10111;
  assign _0680_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:344" *) 5'b11000;
  assign _0681_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:346" *) 5'b11000;
  assign _0682_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:349" *) 5'b11001;
  assign _0683_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) cq_rd9_credits;
  assign _0684_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:351" *) 5'b11001;
  assign _0685_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *) 4'b1001;
  assign _0686_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *) 4'b1000;
  assign _0687_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) 3'b111;
  assign _0688_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) 3'b110;
  assign _0689_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) 3'b101;
  assign _0690_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) 3'b100;
  assign _0691_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) 2'b11;
  assign _0692_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) 2'b10;
  assign _0693_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) 1'b1;
  assign _0694_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3522" *) cq_rd_take_thread_id_last;
  assign _0695_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:354" *) 5'b11010;
  assign _0696_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:356" *) 5'b11010;
  assign _0697_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:359" *) 5'b11011;
  assign _0698_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:361" *) 5'b11011;
  assign _0699_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:364" *) 5'b11100;
  assign _0700_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:366" *) 5'b11100;
  assign _0701_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:369" *) 5'b11101;
  assign _0702_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:371" *) 5'b11101;
  assign _0703_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:374" *) 5'b11110;
  assign _0704_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:376" *) 5'b11110;
  assign _0705_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:379" *) 5'b11111;
  assign _0706_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:381" *) 5'b11111;
  assign _0707_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:384" *) 6'b100000;
  assign _0708_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:386" *) 6'b100000;
  assign _0709_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:389" *) 6'b100001;
  assign _0710_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:391" *) 6'b100001;
  assign _0711_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:394" *) 6'b100010;
  assign _0712_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:396" *) 6'b100010;
  assign _0713_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:399" *) 6'b100011;
  assign _0714_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:401" *) 6'b100011;
  assign _0715_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:404" *) 6'b100100;
  assign _0716_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:406" *) 6'b100100;
  assign _0717_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:409" *) 6'b100101;
  assign _0718_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:411" *) 6'b100101;
  assign _0719_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:414" *) 6'b100110;
  assign _0720_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:416" *) 6'b100110;
  assign _0721_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:419" *) 6'b100111;
  assign _0722_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:421" *) 6'b100111;
  assign _0723_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:424" *) 6'b101000;
  assign _0724_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:426" *) 6'b101000;
  assign _0725_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:429" *) 6'b101001;
  assign _0726_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:431" *) 6'b101001;
  assign _0727_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:434" *) 6'b101010;
  assign _0728_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:436" *) 6'b101010;
  assign _0729_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:439" *) 6'b101011;
  assign _0730_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:441" *) 6'b101011;
  assign _0731_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:444" *) 6'b101100;
  assign _0732_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:446" *) 6'b101100;
  assign _0733_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:449" *) 6'b101101;
  assign _0734_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:451" *) 6'b101101;
  assign _0735_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:454" *) 6'b101110;
  assign _0736_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:456" *) 6'b101110;
  assign _0737_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:459" *) 6'b101111;
  assign _0738_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:461" *) 6'b101111;
  assign _0739_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:464" *) 6'b110000;
  assign _0740_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:466" *) 6'b110000;
  assign _0741_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:469" *) 6'b110001;
  assign _0742_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:471" *) 6'b110001;
  assign _0743_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:474" *) 6'b110010;
  assign _0744_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:476" *) 6'b110010;
  assign _0745_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:479" *) 6'b110011;
  assign _0746_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:481" *) 6'b110011;
  assign _0747_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:484" *) 6'b110100;
  assign _0748_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:486" *) 6'b110100;
  assign _0749_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:489" *) 6'b110101;
  assign _0750_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:491" *) 6'b110101;
  assign _0751_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:494" *) 6'b110110;
  assign _0752_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:496" *) 6'b110110;
  assign _0753_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:499" *) 6'b110111;
  assign _0754_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:501" *) 6'b110111;
  assign _0755_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:504" *) 6'b111000;
  assign _0756_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:506" *) 6'b111000;
  assign _0757_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:509" *) 6'b111001;
  assign _0758_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:511" *) 6'b111001;
  assign _0759_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:514" *) 6'b111010;
  assign _0760_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:516" *) 6'b111010;
  assign _0761_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:519" *) 6'b111011;
  assign _0762_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:521" *) 6'b111011;
  assign _0763_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:524" *) 6'b111100;
  assign _0764_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:526" *) 6'b111100;
  assign _0765_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:529" *) 6'b111101;
  assign _0766_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:531" *) 6'b111101;
  assign _0767_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:534" *) 6'b111110;
  assign _0768_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:536" *) 6'b111110;
  assign _0769_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:539" *) 6'b111111;
  assign _0770_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:541" *) 6'b111111;
  assign _0771_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:544" *) 7'b1000000;
  assign _0772_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:546" *) 7'b1000000;
  assign _0773_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:549" *) 7'b1000001;
  assign _0774_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:551" *) 7'b1000001;
  assign _0775_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:554" *) 7'b1000010;
  assign _0776_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:556" *) 7'b1000010;
  assign _0777_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:559" *) 7'b1000011;
  assign _0778_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:561" *) 7'b1000011;
  assign _0779_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:564" *) 7'b1000100;
  assign _0780_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:566" *) 7'b1000100;
  assign _0781_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:569" *) 7'b1000101;
  assign _0782_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:571" *) 7'b1000101;
  assign _0783_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:574" *) 7'b1000110;
  assign _0784_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:576" *) 7'b1000110;
  assign _0785_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:579" *) 7'b1000111;
  assign _0786_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:581" *) 7'b1000111;
  assign _0787_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:584" *) 7'b1001000;
  assign _0788_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:586" *) 7'b1001000;
  assign _0789_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:589" *) 7'b1001001;
  assign _0790_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:591" *) 7'b1001001;
  assign _0791_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:594" *) 7'b1001010;
  assign _0792_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:596" *) 7'b1001010;
  assign _0793_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:599" *) 7'b1001011;
  assign _0794_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:601" *) 7'b1001011;
  assign _0795_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:604" *) 7'b1001100;
  assign _0796_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:606" *) 7'b1001100;
  assign _0797_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:609" *) 7'b1001101;
  assign _0798_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:611" *) 7'b1001101;
  assign _0799_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:614" *) 7'b1001110;
  assign _0800_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:616" *) 7'b1001110;
  assign _0801_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:619" *) 7'b1001111;
  assign _0802_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:621" *) 7'b1001111;
  assign _0803_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:624" *) 7'b1010000;
  assign _0804_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:626" *) 7'b1010000;
  assign _0805_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:629" *) 7'b1010001;
  assign _0806_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:631" *) 7'b1010001;
  assign _0807_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:634" *) 7'b1010010;
  assign _0808_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:636" *) 7'b1010010;
  assign _0809_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:639" *) 7'b1010011;
  assign _0810_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:641" *) 7'b1010011;
  assign _0811_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:644" *) 7'b1010100;
  assign _0812_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:646" *) 7'b1010100;
  assign _0813_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:649" *) 7'b1010101;
  assign _0814_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:651" *) 7'b1010101;
  assign _0815_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:654" *) 7'b1010110;
  assign _0816_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:656" *) 7'b1010110;
  assign _0817_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:659" *) 7'b1010111;
  assign _0818_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:661" *) 7'b1010111;
  assign _0819_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:664" *) 7'b1011000;
  assign _0820_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:666" *) 7'b1011000;
  assign _0821_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:669" *) 7'b1011001;
  assign _0822_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:671" *) 7'b1011001;
  assign _0823_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:674" *) 7'b1011010;
  assign _0824_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:676" *) 7'b1011010;
  assign _0825_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:679" *) 7'b1011011;
  assign _0826_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:681" *) 7'b1011011;
  assign _0827_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:684" *) 7'b1011100;
  assign _0828_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:686" *) 7'b1011100;
  assign _0829_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:689" *) 7'b1011101;
  assign _0830_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:691" *) 7'b1011101;
  assign _0831_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:694" *) 7'b1011110;
  assign _0832_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:696" *) 7'b1011110;
  assign _0833_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:699" *) 7'b1011111;
  assign _0834_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:701" *) 7'b1011111;
  assign _0835_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:704" *) 7'b1100000;
  assign _0836_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:706" *) 7'b1100000;
  assign _0837_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:709" *) 7'b1100001;
  assign _0838_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:711" *) 7'b1100001;
  assign _0839_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:714" *) 7'b1100010;
  assign _0840_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:716" *) 7'b1100010;
  assign _0841_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:719" *) 7'b1100011;
  assign _0842_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:721" *) 7'b1100011;
  assign _0843_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:724" *) 7'b1100100;
  assign _0844_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:726" *) 7'b1100100;
  assign _0845_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:729" *) 7'b1100101;
  assign _0846_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:731" *) 7'b1100101;
  assign _0847_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:734" *) 7'b1100110;
  assign _0848_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:736" *) 7'b1100110;
  assign _0849_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:739" *) 7'b1100111;
  assign _0850_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:741" *) 7'b1100111;
  assign _0851_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:744" *) 7'b1101000;
  assign _0852_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:746" *) 7'b1101000;
  assign _0853_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:749" *) 7'b1101001;
  assign _0854_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:751" *) 7'b1101001;
  assign _0855_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:754" *) 7'b1101010;
  assign _0856_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:756" *) 7'b1101010;
  assign _0857_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:759" *) 7'b1101011;
  assign _0858_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:761" *) 7'b1101011;
  assign _0859_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:764" *) 7'b1101100;
  assign _0860_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:766" *) 7'b1101100;
  assign _0861_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:769" *) 7'b1101101;
  assign _0862_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:771" *) 7'b1101101;
  assign _0863_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:774" *) 7'b1101110;
  assign _0864_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:776" *) 7'b1101110;
  assign _0865_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:779" *) 7'b1101111;
  assign _0866_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:781" *) 7'b1101111;
  assign _0867_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:784" *) 7'b1110000;
  assign _0868_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:786" *) 7'b1110000;
  assign _0869_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:789" *) 7'b1110001;
  assign _0870_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:791" *) 7'b1110001;
  assign _0871_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:794" *) 7'b1110010;
  assign _0872_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:796" *) 7'b1110010;
  assign _0873_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:799" *) 7'b1110011;
  assign _0874_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:801" *) 7'b1110011;
  assign _0875_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:804" *) 7'b1110100;
  assign _0876_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:806" *) 7'b1110100;
  assign _0877_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:809" *) 7'b1110101;
  assign _0878_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:811" *) 7'b1110101;
  assign _0879_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:814" *) 7'b1110110;
  assign _0880_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:816" *) 7'b1110110;
  assign _0881_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:819" *) 7'b1110111;
  assign _0882_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:821" *) 7'b1110111;
  assign _0883_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:824" *) 7'b1111000;
  assign _0884_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:826" *) 7'b1111000;
  assign _0885_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:829" *) 7'b1111001;
  assign _0886_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:831" *) 7'b1111001;
  assign _0887_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:834" *) 7'b1111010;
  assign _0888_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:836" *) 7'b1111010;
  assign _0889_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:839" *) 7'b1111011;
  assign _0890_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:841" *) 7'b1111011;
  assign _0891_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:844" *) 7'b1111100;
  assign _0892_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:846" *) 7'b1111100;
  assign _0893_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:849" *) 7'b1111101;
  assign _0894_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:851" *) 7'b1111101;
  assign _0895_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:854" *) 7'b1111110;
  assign _0896_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:856" *) 7'b1111110;
  assign _0897_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:859" *) 7'b1111111;
  assign _0898_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:861" *) 7'b1111111;
  assign _0899_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:864" *) 8'b10000000;
  assign _0900_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:866" *) 8'b10000000;
  assign _0901_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:869" *) 8'b10000001;
  assign _0902_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:871" *) 8'b10000001;
  assign _0903_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:874" *) 8'b10000010;
  assign _0904_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:876" *) 8'b10000010;
  assign _0905_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:879" *) 8'b10000011;
  assign _0906_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:881" *) 8'b10000011;
  assign _0907_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:884" *) 8'b10000100;
  assign _0908_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:886" *) 8'b10000100;
  assign _0909_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:889" *) 8'b10000101;
  assign _0910_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:891" *) 8'b10000101;
  assign _0911_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:894" *) 8'b10000110;
  assign _0912_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:896" *) 8'b10000110;
  assign _0913_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:899" *) 8'b10000111;
  assign _0914_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:901" *) 8'b10000111;
  assign _0915_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:904" *) 8'b10001000;
  assign _0916_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:906" *) 8'b10001000;
  assign _0917_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:909" *) 8'b10001001;
  assign _0918_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:911" *) 8'b10001001;
  assign _0919_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:914" *) 8'b10001010;
  assign _0920_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:916" *) 8'b10001010;
  assign _0921_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:919" *) 8'b10001011;
  assign _0922_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:921" *) 8'b10001011;
  assign _0923_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:924" *) 8'b10001100;
  assign _0924_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:926" *) 8'b10001100;
  assign _0925_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:929" *) 8'b10001101;
  assign _0926_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:931" *) 8'b10001101;
  assign _0927_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:934" *) 8'b10001110;
  assign _0928_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:936" *) 8'b10001110;
  assign _0929_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:939" *) 8'b10001111;
  assign _0930_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:941" *) 8'b10001111;
  assign _0931_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:944" *) 8'b10010000;
  assign _0932_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:946" *) 8'b10010000;
  assign _0933_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:949" *) 8'b10010001;
  assign _0934_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:951" *) 8'b10010001;
  assign _0935_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:954" *) 8'b10010010;
  assign _0936_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:956" *) 8'b10010010;
  assign _0937_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:959" *) 8'b10010011;
  assign _0938_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:961" *) 8'b10010011;
  assign _0939_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:964" *) 8'b10010100;
  assign _0940_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:966" *) 8'b10010100;
  assign _0941_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:969" *) 8'b10010101;
  assign _0942_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:971" *) 8'b10010101;
  assign _0943_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:974" *) 8'b10010110;
  assign _0944_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:976" *) 8'b10010110;
  assign _0945_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:979" *) 8'b10010111;
  assign _0946_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:981" *) 8'b10010111;
  assign _0947_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:984" *) 8'b10011000;
  assign _0948_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:986" *) 8'b10011000;
  assign _0949_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:989" *) 8'b10011001;
  assign _0950_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:991" *) 8'b10011001;
  assign _0951_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:994" *) 8'b10011010;
  assign _0952_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:996" *) 8'b10011010;
  assign _0953_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:999" *) 8'b10011011;
  assign _0954_ = cq_rd_count0 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2250" *) 1'b1;
  assign _0955_ = cq_rd_count1 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2251" *) 1'b1;
  assign _0956_ = cq_rd_count2 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2252" *) 1'b1;
  assign _0957_ = cq_rd_count3 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2253" *) 1'b1;
  assign _0958_ = cq_rd_count4 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2254" *) 1'b1;
  assign _0959_ = cq_rd_count5 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2255" *) 1'b1;
  assign _0960_ = cq_rd_count6 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2256" *) 1'b1;
  assign _0961_ = cq_rd_count7 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2257" *) 1'b1;
  assign _0962_ = cq_rd_count8 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2258" *) 1'b1;
  assign _0963_ = cq_rd_count9 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2259" *) 1'b1;
  assign _0964_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1001" *) _0384_;
  assign _0965_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1004" *) _0385_;
  assign _0966_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1006" *) _0386_;
  assign _0967_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1009" *) _0387_;
  assign _0968_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1011" *) _0388_;
  assign _0969_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1014" *) _0389_;
  assign _0970_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1016" *) _0390_;
  assign _0971_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1019" *) _0391_;
  assign _0972_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1021" *) _0392_;
  assign _0973_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1024" *) _0393_;
  assign _0974_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1026" *) _0394_;
  assign _0975_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1029" *) _0395_;
  assign _0976_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1031" *) _0396_;
  assign _0977_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1034" *) _0397_;
  assign _0978_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1036" *) _0398_;
  assign _0979_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1039" *) _0399_;
  assign _0980_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1041" *) _0400_;
  assign _0981_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1044" *) _0401_;
  assign _0982_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1046" *) _0402_;
  assign _0983_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1049" *) _0403_;
  assign _0984_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1051" *) _0404_;
  assign _0985_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1054" *) _0405_;
  assign _0986_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1056" *) _0406_;
  assign _0987_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1059" *) _0407_;
  assign _0988_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1061" *) _0408_;
  assign _0989_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1064" *) _0409_;
  assign _0990_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1066" *) _0410_;
  assign _0991_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1069" *) _0411_;
  assign _0992_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1071" *) _0412_;
  assign _0993_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1074" *) _0413_;
  assign _0994_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1076" *) _0414_;
  assign _0995_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1079" *) _0415_;
  assign _0996_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1081" *) _0416_;
  assign _0997_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1084" *) _0417_;
  assign _0998_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1086" *) _0418_;
  assign _0999_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1089" *) _0419_;
  assign _1000_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1091" *) _0420_;
  assign _1001_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1094" *) _0421_;
  assign _1002_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1096" *) _0422_;
  assign _1003_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1099" *) _0423_;
  assign _1004_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1101" *) _0424_;
  assign _1005_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1104" *) _0425_;
  assign _1006_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1106" *) _0426_;
  assign _1007_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1109" *) _0427_;
  assign _1008_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1111" *) _0428_;
  assign _1009_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1114" *) _0429_;
  assign _1010_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1116" *) _0430_;
  assign _1011_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1119" *) _0431_;
  assign _1012_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1121" *) _0432_;
  assign _1013_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1124" *) _0433_;
  assign _1014_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1126" *) _0434_;
  assign _1015_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1129" *) _0435_;
  assign _1016_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1131" *) _0436_;
  assign _1017_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1134" *) _0437_;
  assign _1018_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1136" *) _0438_;
  assign _1019_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1139" *) _0439_;
  assign _1020_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1141" *) _0440_;
  assign _1021_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1144" *) _0441_;
  assign _1022_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1146" *) _0442_;
  assign _1023_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1149" *) _0443_;
  assign _1024_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1151" *) _0444_;
  assign _1025_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1154" *) _0445_;
  assign _1026_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1156" *) _0446_;
  assign _1027_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1159" *) _0447_;
  assign _1028_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1161" *) _0448_;
  assign _1029_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1164" *) _0449_;
  assign _1030_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1166" *) _0450_;
  assign _1031_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1169" *) _0451_;
  assign _1032_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1171" *) _0452_;
  assign _1033_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1174" *) _0453_;
  assign _1034_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1176" *) _0454_;
  assign _1035_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1179" *) _0455_;
  assign _1036_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1181" *) _0456_;
  assign _1037_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1184" *) _0457_;
  assign _1038_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1186" *) _0458_;
  assign _1039_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1189" *) _0459_;
  assign _1040_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1191" *) _0460_;
  assign _1041_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1194" *) _0461_;
  assign _1042_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1196" *) _0462_;
  assign _1043_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1199" *) _0463_;
  assign _1044_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1201" *) _0464_;
  assign _1045_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1204" *) _0465_;
  assign _1046_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1206" *) _0466_;
  assign _1047_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1209" *) _0467_;
  assign _1048_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1211" *) _0468_;
  assign _1049_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1214" *) _0469_;
  assign _1050_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1216" *) _0470_;
  assign _1051_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1219" *) _0471_;
  assign _1052_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1221" *) _0472_;
  assign _1053_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1224" *) _0473_;
  assign _1054_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1226" *) _0474_;
  assign _1055_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1229" *) _0475_;
  assign _1056_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1231" *) _0476_;
  assign _1057_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1234" *) _0477_;
  assign _1058_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1236" *) _0478_;
  assign _1059_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1239" *) _0479_;
  assign _1060_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1241" *) _0480_;
  assign _1061_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1244" *) _0481_;
  assign _1062_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1246" *) _0482_;
  assign _1063_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1249" *) _0483_;
  assign _1064_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1251" *) _0484_;
  assign _1065_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1254" *) _0485_;
  assign _1066_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1256" *) _0486_;
  assign _1067_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1259" *) _0487_;
  assign _1068_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1261" *) _0488_;
  assign _1069_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1264" *) _0489_;
  assign _1070_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1266" *) _0490_;
  assign _1071_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1269" *) _0491_;
  assign _1072_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1271" *) _0492_;
  assign _1073_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1274" *) _0493_;
  assign _1074_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1276" *) _0494_;
  assign _1075_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1279" *) _0495_;
  assign _1076_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1281" *) _0496_;
  assign _1077_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1284" *) _0497_;
  assign _1078_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1286" *) _0498_;
  assign _1079_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1289" *) _0499_;
  assign _1080_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1291" *) _0500_;
  assign _1081_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1294" *) _0501_;
  assign _1082_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1296" *) _0502_;
  assign _1083_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1299" *) _0503_;
  assign _1084_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1301" *) _0504_;
  assign _1085_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1304" *) _0505_;
  assign _1086_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1306" *) _0506_;
  assign _1087_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1309" *) _0507_;
  assign _1088_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1311" *) _0508_;
  assign _1089_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1314" *) _0509_;
  assign _1090_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1316" *) _0510_;
  assign _1091_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1319" *) _0511_;
  assign _1092_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1321" *) _0512_;
  assign _1093_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1324" *) _0513_;
  assign _1094_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1326" *) _0514_;
  assign _1095_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1329" *) _0515_;
  assign _1096_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1331" *) _0516_;
  assign _1097_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1334" *) _0517_;
  assign _1098_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1336" *) _0518_;
  assign _1099_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1339" *) _0519_;
  assign _1100_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1341" *) _0520_;
  assign _1101_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1344" *) _0521_;
  assign _1102_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1346" *) _0522_;
  assign _1103_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1349" *) _0523_;
  assign _1104_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1351" *) _0524_;
  assign _1105_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1354" *) _0525_;
  assign _1106_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1356" *) _0526_;
  assign _1107_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1359" *) _0527_;
  assign _1108_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1361" *) _0528_;
  assign _1109_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1364" *) _0529_;
  assign _1110_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1366" *) _0530_;
  assign _1111_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1369" *) _0531_;
  assign _1112_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1371" *) _0532_;
  assign _1113_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1374" *) _0533_;
  assign _1114_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1376" *) _0534_;
  assign _1115_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1379" *) _0535_;
  assign _1116_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1381" *) _0536_;
  assign _1117_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1384" *) _0537_;
  assign _1118_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1386" *) _0538_;
  assign _1119_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1389" *) _0539_;
  assign _1120_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1391" *) _0540_;
  assign _1121_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1394" *) _0541_;
  assign _1122_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1396" *) _0542_;
  assign _1123_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1399" *) _0543_;
  assign _1124_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1401" *) _0544_;
  assign _1125_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1404" *) _0545_;
  assign _1126_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1406" *) _0546_;
  assign _1127_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1409" *) _0547_;
  assign _1128_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1411" *) _0548_;
  assign _1129_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1414" *) _0549_;
  assign _1130_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1416" *) _0550_;
  assign _1131_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1419" *) _0551_;
  assign _1132_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1421" *) _0552_;
  assign _1133_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1424" *) _0553_;
  assign _1134_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1426" *) _0554_;
  assign _1135_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1429" *) _0555_;
  assign _1136_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1431" *) _0556_;
  assign _1137_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1434" *) _0557_;
  assign _1138_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1436" *) _0558_;
  assign _1139_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1439" *) _0559_;
  assign _1140_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1441" *) _0560_;
  assign _1141_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1444" *) _0561_;
  assign _1142_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1446" *) _0562_;
  assign _1143_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1449" *) _0563_;
  assign _1144_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1451" *) _0564_;
  assign _1145_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1454" *) _0565_;
  assign _1146_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1456" *) _0566_;
  assign _1147_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1459" *) _0567_;
  assign _1148_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1461" *) _0568_;
  assign _1149_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1464" *) _0569_;
  assign _1150_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1466" *) _0570_;
  assign _1151_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1469" *) _0571_;
  assign _1152_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1471" *) _0572_;
  assign _1153_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1474" *) _0573_;
  assign _1154_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1476" *) _0574_;
  assign _1155_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1479" *) _0575_;
  assign _1156_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1481" *) _0576_;
  assign _1157_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1484" *) _0577_;
  assign _1158_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1486" *) _0578_;
  assign _1159_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1489" *) _0579_;
  assign _1160_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1491" *) _0580_;
  assign _1161_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1494" *) _0581_;
  assign _1162_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1496" *) _0582_;
  assign rd_pushing = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:173" *) _2139_;
  assign rd_pushing0 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2013" *) _0583_;
  assign rd_pushing1 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2014" *) _0584_;
  assign rd_pushing2 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2015" *) _0585_;
  assign rd_pushing3 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2016" *) _0586_;
  assign rd_pushing4 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2017" *) _0587_;
  assign rd_pushing5 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2018" *) _0588_;
  assign rd_pushing6 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2019" *) _0589_;
  assign rd_pushing7 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2020" *) _0590_;
  assign rd_pushing8 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2021" *) _0591_;
  assign rd_pushing9 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2022" *) _0592_;
  assign rd_take0 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2037" *) _0593_;
  assign rd_take1 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2038" *) _0594_;
  assign rd_take2 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2039" *) _0595_;
  assign rd_take3 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2040" *) _0596_;
  assign rd_take4 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2041" *) _0597_;
  assign rd_take5 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2042" *) _0598_;
  assign rd_take6 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2043" *) _0599_;
  assign rd_take7 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2044" *) _0600_;
  assign rd_take8 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2045" *) _0601_;
  assign rd_take9 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2046" *) _0602_;
  assign _1163_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:224" *) _0603_;
  assign update_head_next[0] = rd_take0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2250" *) _0954_;
  assign update_head_next[1] = rd_take1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2251" *) _0955_;
  assign update_head_next[2] = rd_take2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2252" *) _0956_;
  assign update_head_next[3] = rd_take3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2253" *) _0957_;
  assign update_head_next[4] = rd_take4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2254" *) _0958_;
  assign update_head_next[5] = rd_take5 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2255" *) _0959_;
  assign update_head_next[6] = rd_take6 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2256" *) _0960_;
  assign update_head_next[7] = rd_take7 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2257" *) _0961_;
  assign update_head_next[8] = rd_take8 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2258" *) _0962_;
  assign update_head_next[9] = rd_take9 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2259" *) _0963_;
  assign _1164_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:226" *) _0604_;
  assign _1165_ = rd_pushing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2285" *) _0605_;
  assign _1166_ = rd_pushing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *) rd_take0;
  assign _1167_ = _1166_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *) _0606_;
  assign _1168_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:229" *) _0607_;
  assign _1169_ = rd_pushing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2300" *) _0608_;
  assign _1170_ = rd_pushing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *) rd_take1;
  assign _1171_ = _1170_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *) _0609_;
  assign _1172_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:231" *) _0610_;
  assign _1173_ = rd_pushing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2315" *) _0611_;
  assign _1174_ = rd_pushing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *) rd_take2;
  assign _1175_ = _1174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *) _0612_;
  assign _1176_ = rd_pushing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2330" *) _0613_;
  assign _1177_ = rd_pushing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *) rd_take3;
  assign _1178_ = _1177_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *) _0614_;
  assign _1179_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:234" *) _0615_;
  assign _1180_ = rd_pushing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2345" *) _0616_;
  assign _1181_ = rd_pushing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *) rd_take4;
  assign _1182_ = _1181_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *) _0617_;
  assign _1183_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:236" *) _0618_;
  assign _1184_ = rd_pushing5 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2360" *) _0619_;
  assign _1185_ = rd_pushing5 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *) rd_take5;
  assign _1186_ = _1185_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *) _0620_;
  assign _1187_ = rd_pushing6 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2375" *) _0621_;
  assign _1188_ = rd_pushing6 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *) rd_take6;
  assign _1189_ = _1188_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *) _0622_;
  assign _1190_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:239" *) _0623_;
  assign _1191_ = rd_pushing7 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2390" *) _0624_;
  assign _1192_ = rd_pushing7 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *) rd_take7;
  assign _1193_ = _1192_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *) _0625_;
  assign _1194_ = rd_pushing8 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2405" *) _0626_;
  assign _1195_ = rd_pushing8 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *) rd_take8;
  assign _1196_ = _1195_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *) _0627_;
  assign _1197_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:241" *) _0628_;
  assign _1198_ = rd_pushing9 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2420" *) _0629_;
  assign _1199_ = rd_pushing9 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *) rd_take9;
  assign _1200_ = _1199_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *) _0630_;
  assign _1201_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:244" *) _0631_;
  assign _1202_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2457" *) _2447_;
  assign _1203_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2458" *) _2448_;
  assign _1204_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2459" *) _2449_;
  assign _1205_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:246" *) _0632_;
  assign _1206_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2460" *) _2450_;
  assign _1207_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2461" *) _2451_;
  assign _1208_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2462" *) _2452_;
  assign _1209_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2463" *) _2453_;
  assign _1210_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2464" *) _2454_;
  assign _1211_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2465" *) _2455_;
  assign _1212_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2466" *) _2456_;
  assign _1213_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2474" *) _2447_;
  assign _1214_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2475" *) _2448_;
  assign _1215_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2476" *) _2449_;
  assign _1216_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2477" *) _2450_;
  assign _1217_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2478" *) _2451_;
  assign _1218_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2479" *) _2452_;
  assign _1219_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2480" *) _2453_;
  assign _1220_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2481" *) _2454_;
  assign _1221_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2482" *) _2455_;
  assign _1222_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2483" *) _2456_;
  assign _1223_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:249" *) _0633_;
  assign _1224_ = rd_take_n_dly[0] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2491" *) update_head[0];
  assign _1225_ = rd_take_n_dly[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2492" *) update_head[1];
  assign _1226_ = rd_take_n_dly[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2493" *) update_head[2];
  assign _1227_ = rd_take_n_dly[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2494" *) update_head[3];
  assign _1228_ = rd_take_n_dly[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2495" *) update_head[4];
  assign _1229_ = rd_take_n_dly[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2496" *) update_head[5];
  assign _1230_ = rd_take_n_dly[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2497" *) update_head[6];
  assign _1231_ = rd_take_n_dly[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2498" *) update_head[7];
  assign _1232_ = rd_take_n_dly[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2499" *) update_head[8];
  assign _1233_ = rd_take_n_dly[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2500" *) update_head[9];
  assign _1234_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:251" *) _0634_;
  assign _1235_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:254" *) _0635_;
  assign _1236_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:256" *) _0636_;
  assign _1237_ = cq_rd0_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) cq_rd0_prdy;
  assign _1238_ = _1237_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) _2141_;
  assign _1239_ = _2243_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) _2244_;
  assign _1240_ = _1237_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2571" *) rd_skid0_1_vld;
  assign _1241_ = _1237_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *) _2142_;
  assign _1242_ = _2243_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *) _2245_;
  assign _1243_ = _1237_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2583" *) rd_skid0_2_vld;
  assign _1244_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:259" *) _0637_;
  assign _1245_ = _2243_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) rd_skid0_0_vld;
  assign _1246_ = _1245_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) rd_skid0_1_vld;
  assign _1247_ = _1246_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) _2246_;
  assign _1248_ = rd_bypassing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) rd_skid0_0_vld;
  assign _1249_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:261" *) _0638_;
  assign _1250_ = rd_skid0_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *) _2243_;
  assign _1251_ = rd_skid0_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2612" *) _2243_;
  assign _1252_ = _2142_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) _2144_;
  assign cq_rd_take_elig[0] = _2255_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) _2256_;
  assign wr_reserving = cq_wr_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) cq_wr_prdy;
  assign _1253_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) _0583_;
  assign _1254_ = _1253_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) _0639_;
  assign _1255_ = _1254_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) _2145_;
  assign rd_pre_bypassing0 = _1255_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) _2257_;
  assign _1256_ = _2146_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) rd_skid0_0_vld;
  assign _1257_ = _1256_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) rd_skid0_1_vld;
  assign _1258_ = rd_pre_bypassing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) _2259_;
  assign rd_bypassing0 = _1258_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) _2144_;
  assign _1259_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:264" *) _0640_;
  assign _1260_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:266" *) _0641_;
  assign _1261_ = cq_rd1_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) cq_rd1_prdy;
  assign _1262_ = _1261_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) _2149_;
  assign _1263_ = _2260_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) _2261_;
  assign _1264_ = _1261_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2667" *) rd_skid1_1_vld;
  assign _1265_ = _1261_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *) _2150_;
  assign _1266_ = _2260_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *) _2262_;
  assign _1267_ = _1261_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2679" *) rd_skid1_2_vld;
  assign _1268_ = _2260_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) rd_skid1_0_vld;
  assign _1269_ = _1268_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) rd_skid1_1_vld;
  assign _1270_ = _1269_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) _2263_;
  assign _1271_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:269" *) _0642_;
  assign _1272_ = rd_bypassing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) rd_skid1_0_vld;
  assign _1273_ = rd_skid1_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *) _2260_;
  assign _1274_ = rd_skid1_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2708" *) _2260_;
  assign _1275_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:271" *) _0643_;
  assign _1276_ = _2150_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) _2152_;
  assign cq_rd_take_elig[1] = _2272_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) _2273_;
  assign _1277_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) _0584_;
  assign _1278_ = _1277_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) _0644_;
  assign _1279_ = _1278_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) _2153_;
  assign rd_pre_bypassing1 = _1279_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) _2274_;
  assign _1280_ = _2154_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) rd_skid1_0_vld;
  assign _1281_ = _1280_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) rd_skid1_1_vld;
  assign _1282_ = rd_pre_bypassing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) _2276_;
  assign rd_bypassing1 = _1282_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) _2152_;
  assign _1283_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:274" *) _0645_;
  assign _1284_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:276" *) _0646_;
  assign _1285_ = cq_rd2_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) cq_rd2_prdy;
  assign _1286_ = _1285_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) _2157_;
  assign _1287_ = _2277_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) _2278_;
  assign _1288_ = _1285_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2763" *) rd_skid2_1_vld;
  assign _1289_ = _1285_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *) _2158_;
  assign _1290_ = _2277_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *) _2279_;
  assign _1291_ = _1285_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2775" *) rd_skid2_2_vld;
  assign _1292_ = _2277_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) rd_skid2_0_vld;
  assign _1293_ = _1292_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) rd_skid2_1_vld;
  assign _1294_ = _1293_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) _2280_;
  assign _1295_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:279" *) _0647_;
  assign _1296_ = rd_bypassing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) rd_skid2_0_vld;
  assign _1297_ = rd_skid2_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *) _2277_;
  assign _1298_ = rd_skid2_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2804" *) _2277_;
  assign _1299_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:281" *) _0648_;
  assign _1300_ = _2158_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) _2160_;
  assign cq_rd_take_elig[2] = _2289_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) _2290_;
  assign _1301_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) _0585_;
  assign _1302_ = _1301_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) _0649_;
  assign _1303_ = _1302_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) _2161_;
  assign rd_pre_bypassing2 = _1303_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) _2291_;
  assign _1304_ = _2162_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) rd_skid2_0_vld;
  assign _1305_ = _1304_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) rd_skid2_1_vld;
  assign _1306_ = rd_pre_bypassing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) _2293_;
  assign rd_bypassing2 = _1306_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) _2160_;
  assign _1307_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:284" *) _0650_;
  assign _1308_ = cq_rd3_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) cq_rd3_prdy;
  assign _1309_ = _1308_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) _2165_;
  assign _1310_ = _2294_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) _2295_;
  assign _1311_ = _1308_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2859" *) rd_skid3_1_vld;
  assign _1312_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:286" *) _0651_;
  assign _1313_ = _1308_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *) _2166_;
  assign _1314_ = _2294_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *) _2296_;
  assign _1315_ = _1308_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2871" *) rd_skid3_2_vld;
  assign _1316_ = _2294_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) rd_skid3_0_vld;
  assign _1317_ = _1316_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) rd_skid3_1_vld;
  assign _1318_ = _1317_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) _2297_;
  assign _1319_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:289" *) _0652_;
  assign _1320_ = rd_bypassing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) rd_skid3_0_vld;
  assign _1321_ = rd_skid3_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *) _2294_;
  assign _1322_ = rd_skid3_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2900" *) _2294_;
  assign _1323_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:291" *) _0653_;
  assign _1324_ = _2166_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) _2168_;
  assign cq_rd_take_elig[3] = _2306_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) _2307_;
  assign _1325_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) _0586_;
  assign _1326_ = _1325_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) _0654_;
  assign _1327_ = _1326_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) _2169_;
  assign rd_pre_bypassing3 = _1327_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) _2308_;
  assign _1328_ = _2170_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) rd_skid3_0_vld;
  assign _1329_ = _1328_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) rd_skid3_1_vld;
  assign _1330_ = rd_pre_bypassing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) _2310_;
  assign rd_bypassing3 = _1330_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) _2168_;
  assign _1331_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:294" *) _0655_;
  assign _1332_ = cq_rd4_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) cq_rd4_prdy;
  assign _1333_ = _1332_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) _2173_;
  assign _1334_ = _2311_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) _2312_;
  assign _1335_ = _1332_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2955" *) rd_skid4_1_vld;
  assign _1336_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:296" *) _0656_;
  assign _1337_ = _1332_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *) _2174_;
  assign _1338_ = _2311_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *) _2313_;
  assign _1339_ = _1332_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2967" *) rd_skid4_2_vld;
  assign _1340_ = _2311_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) rd_skid4_0_vld;
  assign _1341_ = _1340_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) rd_skid4_1_vld;
  assign _1342_ = _1341_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) _2314_;
  assign _1343_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:299" *) _0657_;
  assign _1344_ = rd_bypassing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) rd_skid4_0_vld;
  assign _1345_ = rd_skid4_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *) _2311_;
  assign _1346_ = rd_skid4_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2996" *) _2311_;
  assign _1347_ = _2174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) _2176_;
  assign cq_rd_take_elig[4] = _2323_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) _2324_;
  assign _1348_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:301" *) _0658_;
  assign _1349_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) _0587_;
  assign _1350_ = _1349_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) _0659_;
  assign _1351_ = _1350_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) _2177_;
  assign rd_pre_bypassing4 = _1351_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) _2325_;
  assign _1352_ = _2178_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) rd_skid4_0_vld;
  assign _1353_ = _1352_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) rd_skid4_1_vld;
  assign _1354_ = rd_pre_bypassing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) _2327_;
  assign rd_bypassing4 = _1354_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) _2176_;
  assign _1355_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:304" *) _0660_;
  assign _1356_ = cq_rd5_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) cq_rd5_prdy;
  assign _1357_ = _1356_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) _2181_;
  assign _1358_ = _2328_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) _2329_;
  assign _1359_ = _1356_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3051" *) rd_skid5_1_vld;
  assign _1360_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:306" *) _0661_;
  assign _1361_ = _1356_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *) _2182_;
  assign _1362_ = _2328_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *) _2330_;
  assign _1363_ = _1356_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3063" *) rd_skid5_2_vld;
  assign _1364_ = _2328_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) rd_skid5_0_vld;
  assign _1365_ = _1364_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) rd_skid5_1_vld;
  assign _1366_ = _1365_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) _2331_;
  assign _1367_ = rd_bypassing5 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) rd_skid5_0_vld;
  assign _1368_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:309" *) _0662_;
  assign _1369_ = rd_skid5_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *) _2328_;
  assign _1370_ = rd_skid5_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3092" *) _2328_;
  assign _1371_ = _2182_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) _2184_;
  assign cq_rd_take_elig[5] = _2340_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) _2341_;
  assign _1372_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) _0588_;
  assign _1373_ = _1372_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) _0663_;
  assign _1374_ = _1373_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) _2185_;
  assign rd_pre_bypassing5 = _1374_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) _2342_;
  assign _1375_ = _2186_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) rd_skid5_0_vld;
  assign _1376_ = _1375_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) rd_skid5_1_vld;
  assign _1377_ = rd_pre_bypassing5 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) _2344_;
  assign rd_bypassing5 = _1377_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) _2184_;
  assign _1378_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:311" *) _0664_;
  assign _1379_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:314" *) _0665_;
  assign _1380_ = cq_rd6_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) cq_rd6_prdy;
  assign _1381_ = _1380_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) _2189_;
  assign _1382_ = _2345_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) _2346_;
  assign _1383_ = _1380_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3147" *) rd_skid6_1_vld;
  assign _1384_ = _1380_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *) _2190_;
  assign _1385_ = _2345_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *) _2347_;
  assign _1386_ = _1380_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3159" *) rd_skid6_2_vld;
  assign _1387_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:316" *) _0666_;
  assign _1388_ = _2345_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) rd_skid6_0_vld;
  assign _1389_ = _1388_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) rd_skid6_1_vld;
  assign _1390_ = _1389_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) _2348_;
  assign _1391_ = rd_bypassing6 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) rd_skid6_0_vld;
  assign _1392_ = rd_skid6_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *) _2345_;
  assign _1393_ = rd_skid6_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3188" *) _2345_;
  assign _1394_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:319" *) _0667_;
  assign _1395_ = _2190_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) _2192_;
  assign cq_rd_take_elig[6] = _2357_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) _2358_;
  assign _1396_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) _0589_;
  assign _1397_ = _1396_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) _0668_;
  assign _1398_ = _1397_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) _2193_;
  assign rd_pre_bypassing6 = _1398_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) _2359_;
  assign _1399_ = _2194_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) rd_skid6_0_vld;
  assign _1400_ = _1399_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) rd_skid6_1_vld;
  assign _1401_ = rd_pre_bypassing6 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) _2361_;
  assign rd_bypassing6 = _1401_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) _2192_;
  assign _1402_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:321" *) _0669_;
  assign _1403_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:324" *) _0670_;
  assign _1404_ = cq_rd7_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) cq_rd7_prdy;
  assign _1405_ = _1404_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) _2197_;
  assign _1406_ = _2362_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) _2363_;
  assign _1407_ = _1404_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3243" *) rd_skid7_1_vld;
  assign _1408_ = _1404_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *) _2198_;
  assign _1409_ = _2362_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *) _2364_;
  assign _1410_ = _1404_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3255" *) rd_skid7_2_vld;
  assign _1411_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:326" *) _0671_;
  assign _1412_ = _2362_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) rd_skid7_0_vld;
  assign _1413_ = _1412_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) rd_skid7_1_vld;
  assign _1414_ = _1413_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) _2365_;
  assign _1415_ = rd_bypassing7 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) rd_skid7_0_vld;
  assign _1416_ = rd_skid7_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *) _2362_;
  assign _1417_ = rd_skid7_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3284" *) _2362_;
  assign _1418_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:329" *) _0672_;
  assign _1419_ = _2198_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) _2200_;
  assign cq_rd_take_elig[7] = _2374_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) _2375_;
  assign _1420_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) _0590_;
  assign _1421_ = _1420_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) _0673_;
  assign _1422_ = _1421_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) _2201_;
  assign rd_pre_bypassing7 = _1422_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) _2376_;
  assign _1423_ = _2202_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) rd_skid7_0_vld;
  assign _1424_ = _1423_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) rd_skid7_1_vld;
  assign _1425_ = rd_pre_bypassing7 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) _2378_;
  assign rd_bypassing7 = _1425_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) _2200_;
  assign _1426_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:331" *) _0674_;
  assign _1427_ = cq_rd8_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) cq_rd8_prdy;
  assign _1428_ = _1427_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) _2205_;
  assign _1429_ = _2379_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) _2380_;
  assign _1430_ = _1427_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3339" *) rd_skid8_1_vld;
  assign _1431_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:334" *) _0675_;
  assign _1432_ = _1427_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *) _2206_;
  assign _1433_ = _2379_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *) _2381_;
  assign _1434_ = _1427_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3351" *) rd_skid8_2_vld;
  assign _1435_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:336" *) _0676_;
  assign _1436_ = _2379_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) rd_skid8_0_vld;
  assign _1437_ = _1436_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) rd_skid8_1_vld;
  assign _1438_ = _1437_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) _2382_;
  assign _1439_ = rd_bypassing8 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) rd_skid8_0_vld;
  assign _1440_ = rd_skid8_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *) _2379_;
  assign _1441_ = rd_skid8_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3380" *) _2379_;
  assign _1442_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:339" *) _0677_;
  assign _1443_ = _2206_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) _2208_;
  assign cq_rd_take_elig[8] = _2391_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) _2392_;
  assign _1444_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) _0591_;
  assign _1445_ = _1444_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) _0678_;
  assign _1446_ = _1445_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) _2209_;
  assign rd_pre_bypassing8 = _1446_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) _2393_;
  assign _1447_ = _2210_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) rd_skid8_0_vld;
  assign _1448_ = _1447_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) rd_skid8_1_vld;
  assign _1449_ = rd_pre_bypassing8 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) _2395_;
  assign rd_bypassing8 = _1449_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) _2208_;
  assign _1450_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:341" *) _0679_;
  assign _1451_ = cq_rd9_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) cq_rd9_prdy;
  assign _1452_ = _1451_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) _2213_;
  assign _1453_ = _2396_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) _2397_;
  assign _1454_ = _1451_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3435" *) rd_skid9_1_vld;
  assign _1455_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:344" *) _0680_;
  assign _1456_ = _1451_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *) _2214_;
  assign _1457_ = _2396_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *) _2398_;
  assign _1458_ = _1451_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3447" *) rd_skid9_2_vld;
  assign _1459_ = _2396_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) rd_skid9_0_vld;
  assign _1460_ = _1459_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) rd_skid9_1_vld;
  assign _1461_ = _1460_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) _2399_;
  assign _1462_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:346" *) _0681_;
  assign _1463_ = rd_bypassing9 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) rd_skid9_0_vld;
  assign _1464_ = rd_skid9_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *) _2396_;
  assign _1465_ = rd_skid9_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3476" *) _2396_;
  assign _1466_ = _2214_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) _2216_;
  assign cq_rd_take_elig[9] = _2408_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) _2409_;
  assign _1467_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:349" *) _0682_;
  assign _1468_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) _0592_;
  assign _1469_ = _1468_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) _0683_;
  assign _1470_ = _1469_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) _2217_;
  assign rd_pre_bypassing9 = _1470_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) _2410_;
  assign _1471_ = _2218_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) rd_skid9_0_vld;
  assign _1472_ = _1471_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) rd_skid9_1_vld;
  assign _1473_ = rd_pre_bypassing9 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) _2412_;
  assign rd_bypassing9 = _1473_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) _2216_;
  assign _1474_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:351" *) _0684_;
  assign _1475_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *) _0685_;
  assign cq_rd_take_thread_id_is_1[9] = _1475_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *) _2220_;
  assign _1476_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *) _0686_;
  assign _1477_ = _1476_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *) _2221_;
  assign cq_rd_take_thread_id_is_1[8] = _1477_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *) _2220_;
  assign _1478_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) _0687_;
  assign _1479_ = _1478_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) _2222_;
  assign _1480_ = _1479_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) _2221_;
  assign cq_rd_take_thread_id_is_1[7] = _1480_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) _2220_;
  assign _1481_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) _0688_;
  assign _1482_ = _1481_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) _2223_;
  assign _1483_ = _1482_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) _2222_;
  assign _1484_ = _1483_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) _2221_;
  assign cq_rd_take_thread_id_is_1[6] = _1484_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) _2220_;
  assign _1485_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _0689_;
  assign _1486_ = _1485_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _2224_;
  assign _1487_ = _1486_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _2223_;
  assign _1488_ = _1487_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _2222_;
  assign _1489_ = _1488_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _2221_;
  assign cq_rd_take_thread_id_is_1[5] = _1489_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) _2220_;
  assign _1490_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _0690_;
  assign _1491_ = _1490_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2225_;
  assign _1492_ = _1491_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2224_;
  assign _1493_ = _1492_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2223_;
  assign _1494_ = _1493_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2222_;
  assign _1495_ = _1494_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2221_;
  assign cq_rd_take_thread_id_is_1[4] = _1495_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) _2220_;
  assign _1496_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _0691_;
  assign _1497_ = _1496_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2226_;
  assign _1498_ = _1497_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2225_;
  assign _1499_ = _1498_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2224_;
  assign _1500_ = _1499_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2223_;
  assign _1501_ = _1500_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2222_;
  assign _1502_ = _1501_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2221_;
  assign cq_rd_take_thread_id_is_1[3] = _1502_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) _2220_;
  assign _1503_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _0692_;
  assign _1504_ = _1503_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2227_;
  assign _1505_ = _1504_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2226_;
  assign _1506_ = _1505_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2225_;
  assign _1507_ = _1506_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2224_;
  assign _1508_ = _1507_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2223_;
  assign _1509_ = _1508_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2222_;
  assign _1510_ = _1509_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2221_;
  assign cq_rd_take_thread_id_is_1[2] = _1510_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) _2220_;
  assign _1511_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _0693_;
  assign _1512_ = _1511_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2228_;
  assign _1513_ = _1512_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2227_;
  assign _1514_ = _1513_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2226_;
  assign _1515_ = _1514_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2225_;
  assign _1516_ = _1515_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2224_;
  assign _1517_ = _1516_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2223_;
  assign _1518_ = _1517_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2222_;
  assign _1519_ = _1518_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2221_;
  assign cq_rd_take_thread_id_is_1[1] = _1519_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) _2220_;
  assign cq_rd_take_thread_id_is_1[0] = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3522" *) _0694_;
  assign _1520_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *) _0685_;
  assign _1521_ = _1520_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *) _2220_;
  assign cq_rd_take_thread_id_is_2[9] = _1521_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *) _2229_;
  assign _1522_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *) _0686_;
  assign _1523_ = _1522_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *) _2221_;
  assign _1524_ = _1523_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *) _2220_;
  assign cq_rd_take_thread_id_is_2[8] = _1524_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3525" *) _2229_;
  assign _1525_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *) _0687_;
  assign _1526_ = _1525_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *) _2222_;
  assign _1527_ = _1526_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *) _2221_;
  assign _1528_ = _1527_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *) _2220_;
  assign cq_rd_take_thread_id_is_2[7] = _1528_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3526" *) _2229_;
  assign _1529_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _0688_;
  assign _1530_ = _1529_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _2223_;
  assign _1531_ = _1530_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _2222_;
  assign _1532_ = _1531_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _2221_;
  assign _1533_ = _1532_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _2220_;
  assign cq_rd_take_thread_id_is_2[6] = _1533_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3527" *) _2229_;
  assign _1534_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _0689_;
  assign _1535_ = _1534_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2224_;
  assign _1536_ = _1535_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2223_;
  assign _1537_ = _1536_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2222_;
  assign _1538_ = _1537_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2221_;
  assign _1539_ = _1538_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2220_;
  assign cq_rd_take_thread_id_is_2[5] = _1539_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3528" *) _2229_;
  assign _1540_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _0690_;
  assign _1541_ = _1540_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2225_;
  assign _1542_ = _1541_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2224_;
  assign _1543_ = _1542_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2223_;
  assign _1544_ = _1543_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2222_;
  assign _1545_ = _1544_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2221_;
  assign _1546_ = _1545_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2220_;
  assign cq_rd_take_thread_id_is_2[4] = _1546_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3529" *) _2229_;
  assign _1547_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _0691_;
  assign _1548_ = _1547_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2226_;
  assign _1549_ = _1548_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2225_;
  assign _1550_ = _1549_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2224_;
  assign _1551_ = _1550_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2223_;
  assign _1552_ = _1551_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2222_;
  assign _1553_ = _1552_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2221_;
  assign _1554_ = _1553_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2220_;
  assign cq_rd_take_thread_id_is_2[3] = _1554_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3530" *) _2229_;
  assign _1555_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _0692_;
  assign _1556_ = _1555_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2227_;
  assign _1557_ = _1556_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2226_;
  assign _1558_ = _1557_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2225_;
  assign _1559_ = _1558_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2224_;
  assign _1560_ = _1559_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2223_;
  assign _1561_ = _1560_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2222_;
  assign _1562_ = _1561_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2221_;
  assign _1563_ = _1562_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2220_;
  assign cq_rd_take_thread_id_is_2[2] = _1563_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3531" *) _2229_;
  assign cq_rd_take_thread_id_is_2[1] = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3532" *) _0693_;
  assign _1564_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3533" *) _0694_;
  assign cq_rd_take_thread_id_is_2[0] = _1564_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3533" *) _2229_;
  assign _1565_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *) _0685_;
  assign _1566_ = _1565_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *) _2220_;
  assign _1567_ = _1566_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *) _2229_;
  assign cq_rd_take_thread_id_is_3[9] = _1567_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3535" *) _2228_;
  assign _1568_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *) _0686_;
  assign _1569_ = _1568_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *) _2221_;
  assign _1570_ = _1569_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *) _2220_;
  assign _1571_ = _1570_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *) _2229_;
  assign cq_rd_take_thread_id_is_3[8] = _1571_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3536" *) _2228_;
  assign _1572_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _0687_;
  assign _1573_ = _1572_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _2222_;
  assign _1574_ = _1573_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _2221_;
  assign _1575_ = _1574_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _2220_;
  assign _1576_ = _1575_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _2229_;
  assign cq_rd_take_thread_id_is_3[7] = _1576_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3537" *) _2228_;
  assign _1577_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _0688_;
  assign _1578_ = _1577_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2223_;
  assign _1579_ = _1578_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2222_;
  assign _1580_ = _1579_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2221_;
  assign _1581_ = _1580_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2220_;
  assign _1582_ = _1581_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2229_;
  assign cq_rd_take_thread_id_is_3[6] = _1582_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3538" *) _2228_;
  assign _1583_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _0689_;
  assign _1584_ = _1583_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2224_;
  assign _1585_ = _1584_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2223_;
  assign _1586_ = _1585_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2222_;
  assign _1587_ = _1586_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2221_;
  assign _1588_ = _1587_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2220_;
  assign _1589_ = _1588_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2229_;
  assign cq_rd_take_thread_id_is_3[5] = _1589_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3539" *) _2228_;
  assign _1590_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:354" *) _0695_;
  assign _1591_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _0690_;
  assign _1592_ = _1591_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2225_;
  assign _1593_ = _1592_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2224_;
  assign _1594_ = _1593_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2223_;
  assign _1595_ = _1594_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2222_;
  assign _1596_ = _1595_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2221_;
  assign _1597_ = _1596_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2220_;
  assign _1598_ = _1597_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2229_;
  assign cq_rd_take_thread_id_is_3[4] = _1598_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3540" *) _2228_;
  assign _1599_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _0691_;
  assign _1600_ = _1599_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2226_;
  assign _1601_ = _1600_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2225_;
  assign _1602_ = _1601_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2224_;
  assign _1603_ = _1602_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2223_;
  assign _1604_ = _1603_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2222_;
  assign _1605_ = _1604_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2221_;
  assign _1606_ = _1605_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2220_;
  assign _1607_ = _1606_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2229_;
  assign cq_rd_take_thread_id_is_3[3] = _1607_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3541" *) _2228_;
  assign cq_rd_take_thread_id_is_3[2] = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3542" *) _0692_;
  assign _1608_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3543" *) _0693_;
  assign cq_rd_take_thread_id_is_3[1] = _1608_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3543" *) _2228_;
  assign _1609_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3544" *) _0694_;
  assign _1610_ = _1609_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3544" *) _2229_;
  assign cq_rd_take_thread_id_is_3[0] = _1610_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3544" *) _2228_;
  assign _1611_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *) _0685_;
  assign _1612_ = _1611_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *) _2220_;
  assign _1613_ = _1612_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *) _2229_;
  assign _1614_ = _1613_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *) _2228_;
  assign cq_rd_take_thread_id_is_4[9] = _1614_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3546" *) _2227_;
  assign _1615_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _0686_;
  assign _1616_ = _1615_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _2221_;
  assign _1617_ = _1616_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _2220_;
  assign _1618_ = _1617_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _2229_;
  assign _1619_ = _1618_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _2228_;
  assign cq_rd_take_thread_id_is_4[8] = _1619_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3547" *) _2227_;
  assign _1620_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _0687_;
  assign _1621_ = _1620_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2222_;
  assign _1622_ = _1621_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2221_;
  assign _1623_ = _1622_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2220_;
  assign _1624_ = _1623_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2229_;
  assign _1625_ = _1624_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2228_;
  assign cq_rd_take_thread_id_is_4[7] = _1625_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3548" *) _2227_;
  assign _1626_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _0688_;
  assign _1627_ = _1626_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2223_;
  assign _1628_ = _1627_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2222_;
  assign _1629_ = _1628_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2221_;
  assign _1630_ = _1629_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2220_;
  assign _1631_ = _1630_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2229_;
  assign _1632_ = _1631_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2228_;
  assign cq_rd_take_thread_id_is_4[6] = _1632_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3549" *) _2227_;
  assign _1633_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _0689_;
  assign _1634_ = _1633_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2224_;
  assign _1635_ = _1634_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2223_;
  assign _1636_ = _1635_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2222_;
  assign _1637_ = _1636_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2221_;
  assign _1638_ = _1637_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2220_;
  assign _1639_ = _1638_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2229_;
  assign _1640_ = _1639_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2228_;
  assign cq_rd_take_thread_id_is_4[5] = _1640_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3550" *) _2227_;
  assign _1641_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _0690_;
  assign _1642_ = _1641_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2225_;
  assign _1643_ = _1642_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2224_;
  assign _1644_ = _1643_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2223_;
  assign _1645_ = _1644_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2222_;
  assign _1646_ = _1645_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2221_;
  assign _1647_ = _1646_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2220_;
  assign _1648_ = _1647_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2229_;
  assign _1649_ = _1648_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2228_;
  assign cq_rd_take_thread_id_is_4[4] = _1649_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3551" *) _2227_;
  assign cq_rd_take_thread_id_is_4[3] = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3552" *) _0691_;
  assign _1650_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3553" *) _0692_;
  assign cq_rd_take_thread_id_is_4[2] = _1650_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3553" *) _2227_;
  assign _1651_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3554" *) _0693_;
  assign _1652_ = _1651_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3554" *) _2228_;
  assign cq_rd_take_thread_id_is_4[1] = _1652_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3554" *) _2227_;
  assign _1653_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *) _0694_;
  assign _1654_ = _1653_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *) _2229_;
  assign _1655_ = _1654_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *) _2228_;
  assign cq_rd_take_thread_id_is_4[0] = _1655_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3555" *) _2227_;
  assign _1656_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _0685_;
  assign _1657_ = _1656_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _2220_;
  assign _1658_ = _1657_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _2229_;
  assign _1659_ = _1658_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _2228_;
  assign _1660_ = _1659_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _2227_;
  assign cq_rd_take_thread_id_is_5[9] = _1660_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3557" *) _2226_;
  assign _1661_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _0686_;
  assign _1662_ = _1661_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2221_;
  assign _1663_ = _1662_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2220_;
  assign _1664_ = _1663_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2229_;
  assign _1665_ = _1664_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2228_;
  assign _1666_ = _1665_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2227_;
  assign cq_rd_take_thread_id_is_5[8] = _1666_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3558" *) _2226_;
  assign _1667_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _0687_;
  assign _1668_ = _1667_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2222_;
  assign _1669_ = _1668_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2221_;
  assign _1670_ = _1669_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2220_;
  assign _1671_ = _1670_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2229_;
  assign _1672_ = _1671_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2228_;
  assign _1673_ = _1672_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2227_;
  assign cq_rd_take_thread_id_is_5[7] = _1673_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3559" *) _2226_;
  assign _1674_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:356" *) _0696_;
  assign _1675_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _0688_;
  assign _1676_ = _1675_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2223_;
  assign _1677_ = _1676_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2222_;
  assign _1678_ = _1677_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2221_;
  assign _1679_ = _1678_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2220_;
  assign _1680_ = _1679_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2229_;
  assign _1681_ = _1680_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2228_;
  assign _1682_ = _1681_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2227_;
  assign cq_rd_take_thread_id_is_5[6] = _1682_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3560" *) _2226_;
  assign _1683_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _0689_;
  assign _1684_ = _1683_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2224_;
  assign _1685_ = _1684_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2223_;
  assign _1686_ = _1685_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2222_;
  assign _1687_ = _1686_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2221_;
  assign _1688_ = _1687_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2220_;
  assign _1689_ = _1688_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2229_;
  assign _1690_ = _1689_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2228_;
  assign _1691_ = _1690_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2227_;
  assign cq_rd_take_thread_id_is_5[5] = _1691_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3561" *) _2226_;
  assign cq_rd_take_thread_id_is_5[4] = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3562" *) _0690_;
  assign _1692_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3563" *) _0691_;
  assign cq_rd_take_thread_id_is_5[3] = _1692_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3563" *) _2226_;
  assign _1693_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3564" *) _0692_;
  assign _1694_ = _1693_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3564" *) _2227_;
  assign cq_rd_take_thread_id_is_5[2] = _1694_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3564" *) _2226_;
  assign _1695_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *) _0693_;
  assign _1696_ = _1695_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *) _2228_;
  assign _1697_ = _1696_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *) _2227_;
  assign cq_rd_take_thread_id_is_5[1] = _1697_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3565" *) _2226_;
  assign _1698_ = cq_rd_take_elig[5] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *) _0694_;
  assign _1699_ = _1698_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *) _2229_;
  assign _1700_ = _1699_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *) _2228_;
  assign _1701_ = _1700_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *) _2227_;
  assign cq_rd_take_thread_id_is_5[0] = _1701_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3566" *) _2226_;
  assign _1702_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _0685_;
  assign _1703_ = _1702_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2220_;
  assign _1704_ = _1703_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2229_;
  assign _1705_ = _1704_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2228_;
  assign _1706_ = _1705_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2227_;
  assign _1707_ = _1706_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2226_;
  assign cq_rd_take_thread_id_is_6[9] = _1707_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3568" *) _2225_;
  assign _1708_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _0686_;
  assign _1709_ = _1708_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2221_;
  assign _1710_ = _1709_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2220_;
  assign _1711_ = _1710_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2229_;
  assign _1712_ = _1711_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2228_;
  assign _1713_ = _1712_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2227_;
  assign _1714_ = _1713_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2226_;
  assign cq_rd_take_thread_id_is_6[8] = _1714_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3569" *) _2225_;
  assign _1715_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _0687_;
  assign _1716_ = _1715_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2222_;
  assign _1717_ = _1716_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2221_;
  assign _1718_ = _1717_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2220_;
  assign _1719_ = _1718_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2229_;
  assign _1720_ = _1719_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2228_;
  assign _1721_ = _1720_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2227_;
  assign _1722_ = _1721_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2226_;
  assign cq_rd_take_thread_id_is_6[7] = _1722_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3570" *) _2225_;
  assign _1723_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _0688_;
  assign _1724_ = _1723_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2223_;
  assign _1725_ = _1724_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2222_;
  assign _1726_ = _1725_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2221_;
  assign _1727_ = _1726_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2220_;
  assign _1728_ = _1727_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2229_;
  assign _1729_ = _1728_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2228_;
  assign _1730_ = _1729_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2227_;
  assign _1731_ = _1730_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2226_;
  assign cq_rd_take_thread_id_is_6[6] = _1731_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3571" *) _2225_;
  assign cq_rd_take_thread_id_is_6[5] = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3572" *) _0689_;
  assign _1732_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3573" *) _0690_;
  assign cq_rd_take_thread_id_is_6[4] = _1732_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3573" *) _2225_;
  assign _1733_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3574" *) _0691_;
  assign _1734_ = _1733_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3574" *) _2226_;
  assign cq_rd_take_thread_id_is_6[3] = _1734_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3574" *) _2225_;
  assign _1735_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *) _0692_;
  assign _1736_ = _1735_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *) _2227_;
  assign _1737_ = _1736_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *) _2226_;
  assign cq_rd_take_thread_id_is_6[2] = _1737_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3575" *) _2225_;
  assign _1738_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *) _0693_;
  assign _1739_ = _1738_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *) _2228_;
  assign _1740_ = _1739_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *) _2227_;
  assign _1741_ = _1740_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *) _2226_;
  assign cq_rd_take_thread_id_is_6[1] = _1741_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3576" *) _2225_;
  assign _1742_ = cq_rd_take_elig[6] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _0694_;
  assign _1743_ = _1742_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _2229_;
  assign _1744_ = _1743_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _2228_;
  assign _1745_ = _1744_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _2227_;
  assign _1746_ = _1745_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _2226_;
  assign cq_rd_take_thread_id_is_6[0] = _1746_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3577" *) _2225_;
  assign _1747_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _0685_;
  assign _1748_ = _1747_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2220_;
  assign _1749_ = _1748_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2229_;
  assign _1750_ = _1749_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2228_;
  assign _1751_ = _1750_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2227_;
  assign _1752_ = _1751_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2226_;
  assign _1753_ = _1752_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2225_;
  assign cq_rd_take_thread_id_is_7[9] = _1753_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3579" *) _2224_;
  assign _1754_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _0686_;
  assign _1755_ = _1754_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2221_;
  assign _1756_ = _1755_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2220_;
  assign _1757_ = _1756_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2229_;
  assign _1758_ = _1757_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2228_;
  assign _1759_ = _1758_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2227_;
  assign _1760_ = _1759_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2226_;
  assign _1761_ = _1760_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2225_;
  assign cq_rd_take_thread_id_is_7[8] = _1761_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3580" *) _2224_;
  assign _1762_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _0687_;
  assign _1763_ = _1762_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2222_;
  assign _1764_ = _1763_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2221_;
  assign _1765_ = _1764_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2220_;
  assign _1766_ = _1765_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2229_;
  assign _1767_ = _1766_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2228_;
  assign _1768_ = _1767_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2227_;
  assign _1769_ = _1768_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2226_;
  assign _1770_ = _1769_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2225_;
  assign cq_rd_take_thread_id_is_7[7] = _1770_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3581" *) _2224_;
  assign cq_rd_take_thread_id_is_7[6] = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3582" *) _0688_;
  assign _1771_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3583" *) _0689_;
  assign cq_rd_take_thread_id_is_7[5] = _1771_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3583" *) _2224_;
  assign _1772_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3584" *) _0690_;
  assign _1773_ = _1772_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3584" *) _2225_;
  assign cq_rd_take_thread_id_is_7[4] = _1773_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3584" *) _2224_;
  assign _1774_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *) _0691_;
  assign _1775_ = _1774_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *) _2226_;
  assign _1776_ = _1775_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *) _2225_;
  assign cq_rd_take_thread_id_is_7[3] = _1776_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3585" *) _2224_;
  assign _1777_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *) _0692_;
  assign _1778_ = _1777_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *) _2227_;
  assign _1779_ = _1778_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *) _2226_;
  assign _1780_ = _1779_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *) _2225_;
  assign cq_rd_take_thread_id_is_7[2] = _1780_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3586" *) _2224_;
  assign _1781_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _0693_;
  assign _1782_ = _1781_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _2228_;
  assign _1783_ = _1782_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _2227_;
  assign _1784_ = _1783_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _2226_;
  assign _1785_ = _1784_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _2225_;
  assign cq_rd_take_thread_id_is_7[1] = _1785_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3587" *) _2224_;
  assign _1786_ = cq_rd_take_elig[7] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _0694_;
  assign _1787_ = _1786_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2229_;
  assign _1788_ = _1787_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2228_;
  assign _1789_ = _1788_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2227_;
  assign _1790_ = _1789_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2226_;
  assign _1791_ = _1790_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2225_;
  assign cq_rd_take_thread_id_is_7[0] = _1791_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3588" *) _2224_;
  assign _1792_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:359" *) _0697_;
  assign _1793_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _0685_;
  assign _1794_ = _1793_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2220_;
  assign _1795_ = _1794_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2229_;
  assign _1796_ = _1795_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2228_;
  assign _1797_ = _1796_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2227_;
  assign _1798_ = _1797_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2226_;
  assign _1799_ = _1798_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2225_;
  assign _1800_ = _1799_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2224_;
  assign cq_rd_take_thread_id_is_8[9] = _1800_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3590" *) _2223_;
  assign _1801_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _0686_;
  assign _1802_ = _1801_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2221_;
  assign _1803_ = _1802_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2220_;
  assign _1804_ = _1803_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2229_;
  assign _1805_ = _1804_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2228_;
  assign _1806_ = _1805_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2227_;
  assign _1807_ = _1806_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2226_;
  assign _1808_ = _1807_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2225_;
  assign _1809_ = _1808_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2224_;
  assign cq_rd_take_thread_id_is_8[8] = _1809_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3591" *) _2223_;
  assign cq_rd_take_thread_id_is_8[7] = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3592" *) _0687_;
  assign _1810_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3593" *) _0688_;
  assign cq_rd_take_thread_id_is_8[6] = _1810_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3593" *) _2223_;
  assign _1811_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3594" *) _0689_;
  assign _1812_ = _1811_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3594" *) _2224_;
  assign cq_rd_take_thread_id_is_8[5] = _1812_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3594" *) _2223_;
  assign _1813_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *) _0690_;
  assign _1814_ = _1813_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *) _2225_;
  assign _1815_ = _1814_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *) _2224_;
  assign cq_rd_take_thread_id_is_8[4] = _1815_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3595" *) _2223_;
  assign _1816_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *) _0691_;
  assign _1817_ = _1816_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *) _2226_;
  assign _1818_ = _1817_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *) _2225_;
  assign _1819_ = _1818_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *) _2224_;
  assign cq_rd_take_thread_id_is_8[3] = _1819_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3596" *) _2223_;
  assign _1820_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _0692_;
  assign _1821_ = _1820_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _2227_;
  assign _1822_ = _1821_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _2226_;
  assign _1823_ = _1822_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _2225_;
  assign _1824_ = _1823_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _2224_;
  assign cq_rd_take_thread_id_is_8[2] = _1824_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3597" *) _2223_;
  assign _1825_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _0693_;
  assign _1826_ = _1825_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2228_;
  assign _1827_ = _1826_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2227_;
  assign _1828_ = _1827_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2226_;
  assign _1829_ = _1828_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2225_;
  assign _1830_ = _1829_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2224_;
  assign cq_rd_take_thread_id_is_8[1] = _1830_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3598" *) _2223_;
  assign _1831_ = cq_rd_take_elig[8] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _0694_;
  assign _1832_ = _1831_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2229_;
  assign _1833_ = _1832_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2228_;
  assign _1834_ = _1833_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2227_;
  assign _1835_ = _1834_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2226_;
  assign _1836_ = _1835_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2225_;
  assign _1837_ = _1836_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2224_;
  assign cq_rd_take_thread_id_is_8[0] = _1837_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3599" *) _2223_;
  assign _1838_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _0685_;
  assign _1839_ = _1838_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2220_;
  assign _1840_ = _1839_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2229_;
  assign _1841_ = _1840_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2228_;
  assign _1842_ = _1841_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2227_;
  assign _1843_ = _1842_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2226_;
  assign _1844_ = _1843_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2225_;
  assign _1845_ = _1844_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2224_;
  assign _1846_ = _1845_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2223_;
  assign cq_rd_take_thread_id_is_9[9] = _1846_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3601" *) _2222_;
  assign cq_rd_take_thread_id_is_9[8] = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3602" *) _0686_;
  assign _1847_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3603" *) _0687_;
  assign cq_rd_take_thread_id_is_9[7] = _1847_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3603" *) _2222_;
  assign _1848_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3604" *) _0688_;
  assign _1849_ = _1848_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3604" *) _2223_;
  assign cq_rd_take_thread_id_is_9[6] = _1849_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3604" *) _2222_;
  assign _1850_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *) _0689_;
  assign _1851_ = _1850_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *) _2224_;
  assign _1852_ = _1851_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *) _2223_;
  assign cq_rd_take_thread_id_is_9[5] = _1852_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3605" *) _2222_;
  assign _1853_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *) _0690_;
  assign _1854_ = _1853_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *) _2225_;
  assign _1855_ = _1854_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *) _2224_;
  assign _1856_ = _1855_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *) _2223_;
  assign cq_rd_take_thread_id_is_9[4] = _1856_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3606" *) _2222_;
  assign _1857_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _0691_;
  assign _1858_ = _1857_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _2226_;
  assign _1859_ = _1858_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _2225_;
  assign _1860_ = _1859_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _2224_;
  assign _1861_ = _1860_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _2223_;
  assign cq_rd_take_thread_id_is_9[3] = _1861_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3607" *) _2222_;
  assign _1862_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _0692_;
  assign _1863_ = _1862_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2227_;
  assign _1864_ = _1863_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2226_;
  assign _1865_ = _1864_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2225_;
  assign _1866_ = _1865_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2224_;
  assign _1867_ = _1866_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2223_;
  assign cq_rd_take_thread_id_is_9[2] = _1867_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3608" *) _2222_;
  assign _1868_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _0693_;
  assign _1869_ = _1868_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2228_;
  assign _1870_ = _1869_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2227_;
  assign _1871_ = _1870_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2226_;
  assign _1872_ = _1871_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2225_;
  assign _1873_ = _1872_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2224_;
  assign _1874_ = _1873_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2223_;
  assign cq_rd_take_thread_id_is_9[1] = _1874_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3609" *) _2222_;
  assign _1875_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:361" *) _0698_;
  assign _1876_ = cq_rd_take_elig[9] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _0694_;
  assign _1877_ = _1876_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2229_;
  assign _1878_ = _1877_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2228_;
  assign _1879_ = _1878_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2227_;
  assign _1880_ = _1879_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2226_;
  assign _1881_ = _1880_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2225_;
  assign _1882_ = _1881_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2224_;
  assign _1883_ = _1882_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2223_;
  assign cq_rd_take_thread_id_is_9[0] = _1883_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3610" *) _2222_;
  assign _1884_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:364" *) _0699_;
  assign _1885_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:366" *) _0700_;
  assign _1886_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:369" *) _0701_;
  assign _1887_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:371" *) _0702_;
  assign _1888_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:374" *) _0703_;
  assign _1889_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:376" *) _0704_;
  assign _1890_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:379" *) _0705_;
  assign _1891_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:381" *) _0706_;
  assign _1892_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:384" *) _0707_;
  assign _1893_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:386" *) _0708_;
  assign _1894_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:389" *) _0709_;
  assign _1895_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:391" *) _0710_;
  assign _1896_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:394" *) _0711_;
  assign _1897_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:396" *) _0712_;
  assign _1898_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:399" *) _0713_;
  assign _1899_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:401" *) _0714_;
  assign _1900_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:404" *) _0715_;
  assign _1901_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:406" *) _0716_;
  assign _1902_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:409" *) _0717_;
  assign _1903_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:411" *) _0718_;
  assign _1904_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:414" *) _0719_;
  assign _1905_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:416" *) _0720_;
  assign _1906_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:419" *) _0721_;
  assign _1907_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:421" *) _0722_;
  assign _1908_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:424" *) _0723_;
  assign _1909_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:426" *) _0724_;
  assign _1910_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:429" *) _0725_;
  assign _1911_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:431" *) _0726_;
  assign _1912_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:434" *) _0727_;
  assign _1913_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:436" *) _0728_;
  assign _1914_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:439" *) _0729_;
  assign _1915_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:441" *) _0730_;
  assign _1916_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:444" *) _0731_;
  assign _1917_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:446" *) _0732_;
  assign _1918_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:449" *) _0733_;
  assign _1919_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:451" *) _0734_;
  assign _1920_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:454" *) _0735_;
  assign _1921_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:456" *) _0736_;
  assign _1922_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:459" *) _0737_;
  assign _1923_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:461" *) _0738_;
  assign _1924_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:464" *) _0739_;
  assign _1925_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:466" *) _0740_;
  assign _1926_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:469" *) _0741_;
  assign _1927_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:471" *) _0742_;
  assign _1928_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:474" *) _0743_;
  assign _1929_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:476" *) _0744_;
  assign _1930_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:479" *) _0745_;
  assign _1931_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:481" *) _0746_;
  assign _1932_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:484" *) _0747_;
  assign _1933_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:486" *) _0748_;
  assign _1934_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:489" *) _0749_;
  assign _1935_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:491" *) _0750_;
  assign _1936_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:494" *) _0751_;
  assign _1937_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:496" *) _0752_;
  assign _1938_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:499" *) _0753_;
  assign _1939_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:501" *) _0754_;
  assign _1940_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:504" *) _0755_;
  assign _1941_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:506" *) _0756_;
  assign _1942_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:509" *) _0757_;
  assign _1943_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:511" *) _0758_;
  assign _1944_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:514" *) _0759_;
  assign _1945_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:516" *) _0760_;
  assign _1946_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:519" *) _0761_;
  assign _1947_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:521" *) _0762_;
  assign _1948_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:524" *) _0763_;
  assign _1949_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:526" *) _0764_;
  assign _1950_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:529" *) _0765_;
  assign _1951_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:531" *) _0766_;
  assign _1952_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:534" *) _0767_;
  assign _1953_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:536" *) _0768_;
  assign _1954_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:539" *) _0769_;
  assign _1955_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:541" *) _0770_;
  assign _1956_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:544" *) _0771_;
  assign _1957_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:546" *) _0772_;
  assign _1958_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:549" *) _0773_;
  assign _1959_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:551" *) _0774_;
  assign _1960_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:554" *) _0775_;
  assign _1961_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:556" *) _0776_;
  assign _1962_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:559" *) _0777_;
  assign _1963_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:561" *) _0778_;
  assign _1964_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:564" *) _0779_;
  assign _1965_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:566" *) _0780_;
  assign _1966_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:569" *) _0781_;
  assign _1967_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:571" *) _0782_;
  assign _1968_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:574" *) _0783_;
  assign _1969_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:576" *) _0784_;
  assign _1970_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:579" *) _0785_;
  assign _1971_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:581" *) _0786_;
  assign _1972_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:584" *) _0787_;
  assign _1973_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:586" *) _0788_;
  assign _1974_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:589" *) _0789_;
  assign _1975_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:591" *) _0790_;
  assign _1976_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:594" *) _0791_;
  assign _1977_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:596" *) _0792_;
  assign _1978_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:599" *) _0793_;
  assign _1979_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:601" *) _0794_;
  assign _1980_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:604" *) _0795_;
  assign _1981_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:606" *) _0796_;
  assign _1982_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:609" *) _0797_;
  assign _1983_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:611" *) _0798_;
  assign _1984_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:614" *) _0799_;
  assign _1985_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:616" *) _0800_;
  assign _1986_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:619" *) _0801_;
  assign _1987_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:621" *) _0802_;
  assign _1988_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:624" *) _0803_;
  assign _1989_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:626" *) _0804_;
  assign _1990_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:629" *) _0805_;
  assign _1991_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:631" *) _0806_;
  assign _1992_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:634" *) _0807_;
  assign _1993_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:636" *) _0808_;
  assign _1994_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:639" *) _0809_;
  assign _1995_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:641" *) _0810_;
  assign _1996_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:644" *) _0811_;
  assign _1997_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:646" *) _0812_;
  assign _1998_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:649" *) _0813_;
  assign _1999_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:651" *) _0814_;
  assign _2000_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:654" *) _0815_;
  assign _2001_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:656" *) _0816_;
  assign _2002_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:659" *) _0817_;
  assign _2003_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:661" *) _0818_;
  assign _2004_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:664" *) _0819_;
  assign _2005_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:666" *) _0820_;
  assign _2006_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:669" *) _0821_;
  assign _2007_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:671" *) _0822_;
  assign _2008_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:674" *) _0823_;
  assign _2009_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:676" *) _0824_;
  assign _2010_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:679" *) _0825_;
  assign _2011_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:681" *) _0826_;
  assign _2012_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:684" *) _0827_;
  assign _2013_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:686" *) _0828_;
  assign _2014_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:689" *) _0829_;
  assign _2015_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:691" *) _0830_;
  assign _2016_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:694" *) _0831_;
  assign _2017_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:696" *) _0832_;
  assign _2018_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:699" *) _0833_;
  assign _2019_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:701" *) _0834_;
  assign _2020_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:704" *) _0835_;
  assign _2021_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:706" *) _0836_;
  assign _2022_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:709" *) _0837_;
  assign _2023_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:711" *) _0838_;
  assign _2024_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:714" *) _0839_;
  assign _2025_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:716" *) _0840_;
  assign _2026_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:719" *) _0841_;
  assign _2027_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:721" *) _0842_;
  assign _2028_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:724" *) _0843_;
  assign _2029_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:726" *) _0844_;
  assign _2030_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:729" *) _0845_;
  assign _2031_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:731" *) _0846_;
  assign _2032_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:734" *) _0847_;
  assign _2033_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:736" *) _0848_;
  assign _2034_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:739" *) _0849_;
  assign _2035_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:741" *) _0850_;
  assign _2036_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:744" *) _0851_;
  assign _2037_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:746" *) _0852_;
  assign _2038_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:749" *) _0853_;
  assign _2039_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:751" *) _0854_;
  assign _2040_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:754" *) _0855_;
  assign _2041_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:756" *) _0856_;
  assign _2042_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:759" *) _0857_;
  assign _2043_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:761" *) _0858_;
  assign _2044_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:764" *) _0859_;
  assign _2045_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:766" *) _0860_;
  assign _2046_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:769" *) _0861_;
  assign _2047_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:771" *) _0862_;
  assign _2048_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:774" *) _0863_;
  assign _2049_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:776" *) _0864_;
  assign _2050_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:779" *) _0865_;
  assign _2051_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:781" *) _0866_;
  assign _2052_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:784" *) _0867_;
  assign _2053_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:786" *) _0868_;
  assign _2054_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:789" *) _0869_;
  assign _2055_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:791" *) _0870_;
  assign _2056_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:794" *) _0871_;
  assign _2057_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:796" *) _0872_;
  assign _2058_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:799" *) _0873_;
  assign _2059_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:801" *) _0874_;
  assign _2060_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:804" *) _0875_;
  assign _2061_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:806" *) _0876_;
  assign _2062_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:809" *) _0877_;
  assign _2063_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:811" *) _0878_;
  assign _2064_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:814" *) _0879_;
  assign _2065_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:816" *) _0880_;
  assign _2066_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:819" *) _0881_;
  assign _2067_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:821" *) _0882_;
  assign _2068_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:824" *) _0883_;
  assign _2069_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:826" *) _0884_;
  assign _2070_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:829" *) _0885_;
  assign _2071_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:831" *) _0886_;
  assign _2072_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:834" *) _0887_;
  assign _2073_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:836" *) _0888_;
  assign _2074_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:839" *) _0889_;
  assign _2075_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:841" *) _0890_;
  assign _2076_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:844" *) _0891_;
  assign _2077_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:846" *) _0892_;
  assign _2078_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:849" *) _0893_;
  assign _2079_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:851" *) _0894_;
  assign _2080_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:854" *) _0895_;
  assign _2081_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:856" *) _0896_;
  assign _2082_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:859" *) _0897_;
  assign _2083_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:861" *) _0898_;
  assign _2084_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:864" *) _0899_;
  assign _2085_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:866" *) _0900_;
  assign _2086_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:869" *) _0901_;
  assign _2087_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:871" *) _0902_;
  assign _2088_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:874" *) _0903_;
  assign _2089_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:876" *) _0904_;
  assign _2090_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:879" *) _0905_;
  assign _2091_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:881" *) _0906_;
  assign _2092_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:884" *) _0907_;
  assign _2093_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:886" *) _0908_;
  assign _2094_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:889" *) _0909_;
  assign _2095_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:891" *) _0910_;
  assign _2096_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:894" *) _0911_;
  assign _2097_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:896" *) _0912_;
  assign _2098_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:899" *) _0913_;
  assign _2099_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:901" *) _0914_;
  assign _2100_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:904" *) _0915_;
  assign _2101_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:906" *) _0916_;
  assign _2102_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:909" *) _0917_;
  assign _2103_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:911" *) _0918_;
  assign _2104_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:914" *) _0919_;
  assign _2105_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:916" *) _0920_;
  assign _2106_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:919" *) _0921_;
  assign _2107_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:921" *) _0922_;
  assign _2108_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:924" *) _0923_;
  assign _2109_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:926" *) _0924_;
  assign _2110_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:929" *) _0925_;
  assign _2111_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:931" *) _0926_;
  assign _2112_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:934" *) _0927_;
  assign _2113_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:936" *) _0928_;
  assign _2114_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:939" *) _0929_;
  assign _2115_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:941" *) _0930_;
  assign _2116_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:944" *) _0931_;
  assign _2117_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:946" *) _0932_;
  assign _2118_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:949" *) _0933_;
  assign _2119_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:951" *) _0934_;
  assign _2120_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:954" *) _0935_;
  assign _2121_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:956" *) _0936_;
  assign _2122_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:959" *) _0937_;
  assign _2123_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:961" *) _0938_;
  assign _2124_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:964" *) _0939_;
  assign _2125_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:966" *) _0940_;
  assign _2126_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:969" *) _0941_;
  assign _2127_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:971" *) _0942_;
  assign _2128_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:974" *) _0943_;
  assign _2129_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:976" *) _0944_;
  assign _2130_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:979" *) _0945_;
  assign _2131_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:981" *) _0946_;
  assign _2132_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:984" *) _0947_;
  assign _2133_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:986" *) _0948_;
  assign _2134_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:989" *) _0949_;
  assign _2135_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:991" *) _0950_;
  assign _2136_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:994" *) _0951_;
  assign _2137_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:996" *) _0952_;
  assign _2138_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:999" *) _0953_;
  assign cq_wr_prdy = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:121" *) cq_wr_busy_int;
  assign _2139_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:125" *) wr_bypassing;
  assign index_l0_0 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1747" *) free_adr_mask[0];
  assign index_l0_1 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1748" *) free_adr_mask[2];
  assign index_l0_2 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1749" *) free_adr_mask[4];
  assign index_l0_3 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1750" *) free_adr_mask[6];
  assign index_l0_4 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1751" *) free_adr_mask[8];
  assign index_l0_5 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1752" *) free_adr_mask[10];
  assign index_l0_6 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1753" *) free_adr_mask[12];
  assign index_l0_7 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1754" *) free_adr_mask[14];
  assign index_l0_8 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1755" *) free_adr_mask[16];
  assign index_l0_9 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1756" *) free_adr_mask[18];
  assign index_l0_10 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1757" *) free_adr_mask[20];
  assign index_l0_11 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1758" *) free_adr_mask[22];
  assign index_l0_12 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1759" *) free_adr_mask[24];
  assign index_l0_13 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1760" *) free_adr_mask[26];
  assign index_l0_14 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1761" *) free_adr_mask[28];
  assign index_l0_15 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1762" *) free_adr_mask[30];
  assign index_l0_16 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1763" *) free_adr_mask[32];
  assign index_l0_17 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1764" *) free_adr_mask[34];
  assign index_l0_18 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1765" *) free_adr_mask[36];
  assign index_l0_19 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1766" *) free_adr_mask[38];
  assign index_l0_20 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1767" *) free_adr_mask[40];
  assign index_l0_21 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1768" *) free_adr_mask[42];
  assign index_l0_22 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1769" *) free_adr_mask[44];
  assign index_l0_23 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1770" *) free_adr_mask[46];
  assign index_l0_24 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1771" *) free_adr_mask[48];
  assign index_l0_25 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1772" *) free_adr_mask[50];
  assign index_l0_26 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1773" *) free_adr_mask[52];
  assign index_l0_27 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1774" *) free_adr_mask[54];
  assign index_l0_28 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1775" *) free_adr_mask[56];
  assign index_l0_29 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1776" *) free_adr_mask[58];
  assign index_l0_30 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1777" *) free_adr_mask[60];
  assign index_l0_31 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1778" *) free_adr_mask[62];
  assign index_l0_32 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1779" *) free_adr_mask[64];
  assign index_l0_33 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1780" *) free_adr_mask[66];
  assign index_l0_34 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1781" *) free_adr_mask[68];
  assign index_l0_35 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1782" *) free_adr_mask[70];
  assign index_l0_36 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1783" *) free_adr_mask[72];
  assign index_l0_37 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1784" *) free_adr_mask[74];
  assign index_l0_38 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1785" *) free_adr_mask[76];
  assign index_l0_39 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1786" *) free_adr_mask[78];
  assign index_l0_40 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1787" *) free_adr_mask[80];
  assign index_l0_41 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1788" *) free_adr_mask[82];
  assign index_l0_42 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1789" *) free_adr_mask[84];
  assign index_l0_43 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1790" *) free_adr_mask[86];
  assign index_l0_44 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1791" *) free_adr_mask[88];
  assign index_l0_45 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1792" *) free_adr_mask[90];
  assign index_l0_46 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1793" *) free_adr_mask[92];
  assign index_l0_47 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1794" *) free_adr_mask[94];
  assign index_l0_48 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1795" *) free_adr_mask[96];
  assign index_l0_49 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1796" *) free_adr_mask[98];
  assign index_l0_50 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1797" *) free_adr_mask[100];
  assign index_l0_51 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1798" *) free_adr_mask[102];
  assign index_l0_52 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1799" *) free_adr_mask[104];
  assign index_l0_53 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1800" *) free_adr_mask[106];
  assign index_l0_54 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1801" *) free_adr_mask[108];
  assign index_l0_55 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1802" *) free_adr_mask[110];
  assign index_l0_56 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1803" *) free_adr_mask[112];
  assign index_l0_57 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1804" *) free_adr_mask[114];
  assign index_l0_58 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1805" *) free_adr_mask[116];
  assign index_l0_59 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1806" *) free_adr_mask[118];
  assign index_l0_60 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1807" *) free_adr_mask[120];
  assign index_l0_61 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1808" *) free_adr_mask[122];
  assign index_l0_62 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1809" *) free_adr_mask[124];
  assign index_l0_63 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1810" *) free_adr_mask[126];
  assign index_l0_64 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1811" *) free_adr_mask[128];
  assign index_l0_65 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1812" *) free_adr_mask[130];
  assign index_l0_66 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1813" *) free_adr_mask[132];
  assign index_l0_67 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1814" *) free_adr_mask[134];
  assign index_l0_68 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1815" *) free_adr_mask[136];
  assign index_l0_69 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1816" *) free_adr_mask[138];
  assign index_l0_70 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1817" *) free_adr_mask[140];
  assign index_l0_71 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1818" *) free_adr_mask[142];
  assign index_l0_72 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1819" *) free_adr_mask[144];
  assign index_l0_73 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1820" *) free_adr_mask[146];
  assign index_l0_74 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1821" *) free_adr_mask[148];
  assign index_l0_75 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1822" *) free_adr_mask[150];
  assign index_l0_76 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1823" *) free_adr_mask[152];
  assign index_l0_77 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1824" *) free_adr_mask[154];
  assign index_l0_78 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1825" *) free_adr_mask[156];
  assign index_l0_79 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1826" *) free_adr_mask[158];
  assign index_l0_80 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1827" *) free_adr_mask[160];
  assign index_l0_81 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1828" *) free_adr_mask[162];
  assign index_l0_82 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1829" *) free_adr_mask[164];
  assign index_l0_83 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1830" *) free_adr_mask[166];
  assign index_l0_84 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1831" *) free_adr_mask[168];
  assign index_l0_85 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1832" *) free_adr_mask[170];
  assign index_l0_86 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1833" *) free_adr_mask[172];
  assign index_l0_87 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1834" *) free_adr_mask[174];
  assign index_l0_88 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1835" *) free_adr_mask[176];
  assign index_l0_89 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1836" *) free_adr_mask[178];
  assign index_l0_90 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1837" *) free_adr_mask[180];
  assign index_l0_91 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1838" *) free_adr_mask[182];
  assign index_l0_92 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1839" *) free_adr_mask[184];
  assign index_l0_93 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1840" *) free_adr_mask[186];
  assign index_l0_94 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1841" *) free_adr_mask[188];
  assign index_l0_95 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1842" *) free_adr_mask[190];
  assign index_l0_96 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1843" *) free_adr_mask[192];
  assign index_l0_97 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1844" *) free_adr_mask[194];
  assign index_l0_98 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1845" *) free_adr_mask[196];
  assign index_l0_99 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1846" *) free_adr_mask[198];
  assign index_l0_100 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1847" *) free_adr_mask[200];
  assign index_l0_101 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1848" *) free_adr_mask[202];
  assign index_l0_102 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1849" *) free_adr_mask[204];
  assign index_l0_103 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1850" *) free_adr_mask[206];
  assign index_l0_104 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1851" *) free_adr_mask[208];
  assign index_l0_105 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1852" *) free_adr_mask[210];
  assign index_l0_106 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1853" *) free_adr_mask[212];
  assign index_l0_107 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1854" *) free_adr_mask[214];
  assign index_l0_108 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1855" *) free_adr_mask[216];
  assign index_l0_109 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1856" *) free_adr_mask[218];
  assign index_l0_110 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1857" *) free_adr_mask[220];
  assign index_l0_111 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1858" *) free_adr_mask[222];
  assign index_l0_112 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1859" *) free_adr_mask[224];
  assign index_l0_113 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1860" *) free_adr_mask[226];
  assign index_l0_114 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1861" *) free_adr_mask[228];
  assign index_l0_115 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1862" *) free_adr_mask[230];
  assign index_l0_116 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1863" *) free_adr_mask[232];
  assign index_l0_117 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1864" *) free_adr_mask[234];
  assign index_l0_118 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1865" *) free_adr_mask[236];
  assign index_l0_119 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1866" *) free_adr_mask[238];
  assign index_l0_120 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1867" *) free_adr_mask[240];
  assign index_l0_121 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1868" *) free_adr_mask[242];
  assign index_l0_122 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1869" *) free_adr_mask[244];
  assign index_l0_123 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1870" *) free_adr_mask[246];
  assign index_l0_124 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1871" *) free_adr_mask[248];
  assign index_l0_125 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1872" *) free_adr_mask[250];
  assign index_l0_126 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1873" *) free_adr_mask[252];
  assign index_l0_127 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1874" *) free_adr_mask[254];
  assign index_l1_0[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1875" *) flag_l0_0;
  assign index_l1_1[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1876" *) flag_l0_2;
  assign index_l1_2[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1877" *) flag_l0_4;
  assign index_l1_3[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1878" *) flag_l0_6;
  assign index_l1_4[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1879" *) flag_l0_8;
  assign index_l1_5[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1880" *) flag_l0_10;
  assign index_l1_6[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1881" *) flag_l0_12;
  assign index_l1_7[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1882" *) flag_l0_14;
  assign index_l1_8[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1883" *) flag_l0_16;
  assign index_l1_9[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1884" *) flag_l0_18;
  assign index_l1_10[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1885" *) flag_l0_20;
  assign index_l1_11[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1886" *) flag_l0_22;
  assign index_l1_12[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1887" *) flag_l0_24;
  assign index_l1_13[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1888" *) flag_l0_26;
  assign index_l1_14[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1889" *) flag_l0_28;
  assign index_l1_15[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1890" *) flag_l0_30;
  assign index_l1_16[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1891" *) flag_l0_32;
  assign index_l1_17[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1892" *) flag_l0_34;
  assign index_l1_18[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1893" *) flag_l0_36;
  assign index_l1_19[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1894" *) flag_l0_38;
  assign index_l1_20[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1895" *) flag_l0_40;
  assign index_l1_21[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1896" *) flag_l0_42;
  assign index_l1_22[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1897" *) flag_l0_44;
  assign index_l1_23[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1898" *) flag_l0_46;
  assign index_l1_24[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1899" *) flag_l0_48;
  assign index_l1_25[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1900" *) flag_l0_50;
  assign index_l1_26[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1901" *) flag_l0_52;
  assign index_l1_27[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1902" *) flag_l0_54;
  assign index_l1_28[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1903" *) flag_l0_56;
  assign index_l1_29[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1904" *) flag_l0_58;
  assign index_l1_30[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1905" *) flag_l0_60;
  assign index_l1_31[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1906" *) flag_l0_62;
  assign index_l1_32[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1907" *) flag_l0_64;
  assign index_l1_33[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1908" *) flag_l0_66;
  assign index_l1_34[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1909" *) flag_l0_68;
  assign index_l1_35[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1910" *) flag_l0_70;
  assign index_l1_36[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1911" *) flag_l0_72;
  assign index_l1_37[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1912" *) flag_l0_74;
  assign index_l1_38[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1913" *) flag_l0_76;
  assign index_l1_39[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1914" *) flag_l0_78;
  assign index_l1_40[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1915" *) flag_l0_80;
  assign index_l1_41[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1916" *) flag_l0_82;
  assign index_l1_42[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1917" *) flag_l0_84;
  assign index_l1_43[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1918" *) flag_l0_86;
  assign index_l1_44[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1919" *) flag_l0_88;
  assign index_l1_45[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1920" *) flag_l0_90;
  assign index_l1_46[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1921" *) flag_l0_92;
  assign index_l1_47[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1922" *) flag_l0_94;
  assign index_l1_48[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1923" *) flag_l0_96;
  assign index_l1_49[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1924" *) flag_l0_98;
  assign index_l1_50[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1925" *) flag_l0_100;
  assign index_l1_51[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1926" *) flag_l0_102;
  assign index_l1_52[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1927" *) flag_l0_104;
  assign index_l1_53[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1928" *) flag_l0_106;
  assign index_l1_54[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1929" *) flag_l0_108;
  assign index_l1_55[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1930" *) flag_l0_110;
  assign index_l1_56[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1931" *) flag_l0_112;
  assign index_l1_57[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1932" *) flag_l0_114;
  assign index_l1_58[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1933" *) flag_l0_116;
  assign index_l1_59[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1934" *) flag_l0_118;
  assign index_l1_60[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1935" *) flag_l0_120;
  assign index_l1_61[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1936" *) flag_l0_122;
  assign index_l1_62[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1937" *) flag_l0_124;
  assign index_l1_63[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1938" *) flag_l0_126;
  assign index_l2_0[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1939" *) flag_l1_0;
  assign index_l2_1[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1940" *) flag_l1_2;
  assign index_l2_2[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1941" *) flag_l1_4;
  assign index_l2_3[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1942" *) flag_l1_6;
  assign index_l2_4[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1943" *) flag_l1_8;
  assign index_l2_5[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1944" *) flag_l1_10;
  assign index_l2_6[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1945" *) flag_l1_12;
  assign index_l2_7[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1946" *) flag_l1_14;
  assign index_l2_8[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1947" *) flag_l1_16;
  assign index_l2_9[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1948" *) flag_l1_18;
  assign index_l2_10[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1949" *) flag_l1_20;
  assign index_l2_11[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1950" *) flag_l1_22;
  assign index_l2_12[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1951" *) flag_l1_24;
  assign index_l2_13[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1952" *) flag_l1_26;
  assign index_l2_14[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1953" *) flag_l1_28;
  assign index_l2_15[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1954" *) flag_l1_30;
  assign index_l2_16[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1955" *) flag_l1_32;
  assign index_l2_17[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1956" *) flag_l1_34;
  assign index_l2_18[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1957" *) flag_l1_36;
  assign index_l2_19[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1958" *) flag_l1_38;
  assign index_l2_20[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1959" *) flag_l1_40;
  assign index_l2_21[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1960" *) flag_l1_42;
  assign index_l2_22[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1961" *) flag_l1_44;
  assign index_l2_23[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1962" *) flag_l1_46;
  assign index_l2_24[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1963" *) flag_l1_48;
  assign index_l2_25[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1964" *) flag_l1_50;
  assign index_l2_26[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1965" *) flag_l1_52;
  assign index_l2_27[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1966" *) flag_l1_54;
  assign index_l2_28[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1967" *) flag_l1_56;
  assign index_l2_29[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1968" *) flag_l1_58;
  assign index_l2_30[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1969" *) flag_l1_60;
  assign index_l2_31[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1970" *) flag_l1_62;
  assign index_l3_0[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1971" *) flag_l2_0;
  assign index_l3_1[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1972" *) flag_l2_2;
  assign index_l3_2[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1973" *) flag_l2_4;
  assign index_l3_3[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1974" *) flag_l2_6;
  assign index_l3_4[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1975" *) flag_l2_8;
  assign index_l3_5[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1976" *) flag_l2_10;
  assign index_l3_6[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1977" *) flag_l2_12;
  assign index_l3_7[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1978" *) flag_l2_14;
  assign index_l3_8[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1979" *) flag_l2_16;
  assign index_l3_9[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1980" *) flag_l2_18;
  assign index_l3_10[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1981" *) flag_l2_20;
  assign index_l3_11[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1982" *) flag_l2_22;
  assign index_l3_12[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1983" *) flag_l2_24;
  assign index_l3_13[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1984" *) flag_l2_26;
  assign index_l3_14[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1985" *) flag_l2_28;
  assign index_l3_15[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1986" *) flag_l2_30;
  assign index_l4_0[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1987" *) flag_l3_0;
  assign index_l4_1[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1988" *) flag_l3_2;
  assign index_l4_2[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1989" *) flag_l3_4;
  assign index_l4_3[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1990" *) flag_l3_6;
  assign index_l4_4[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1991" *) flag_l3_8;
  assign index_l4_5[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1992" *) flag_l3_10;
  assign index_l4_6[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1993" *) flag_l3_12;
  assign index_l4_7[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1994" *) flag_l3_14;
  assign index_l5_0[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1995" *) flag_l4_0;
  assign index_l5_1[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1996" *) flag_l4_2;
  assign index_l5_2[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1997" *) flag_l4_4;
  assign index_l5_3[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1998" *) flag_l4_6;
  assign index_l6_0[6] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1999" *) flag_l5_0;
  assign index_l6_1[6] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2000" *) flag_l5_2;
  assign adr_ram_wr_data[7] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2001" *) flag_l6_0;
  assign _2140_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) rd_skid0_0_vld;
  assign _2141_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) rd_skid0_1_vld;
  assign _2142_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *) rd_skid0_2_vld;
  assign _2143_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) _1237_;
  assign _2144_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) rd_take_n_dly[0];
  assign _2145_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) cq_rd_credit[0];
  assign _2146_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) cq_rd0_prdy_d;
  assign _2147_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) _1257_;
  assign _2148_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) rd_skid1_0_vld;
  assign _2149_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) rd_skid1_1_vld;
  assign _2150_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *) rd_skid1_2_vld;
  assign _2151_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) _1261_;
  assign _2152_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) rd_take_n_dly[1];
  assign _2153_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) cq_rd_credit[1];
  assign _2154_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) cq_rd1_prdy_d;
  assign _2155_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) _1281_;
  assign _2156_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) rd_skid2_0_vld;
  assign _2157_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) rd_skid2_1_vld;
  assign _2158_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *) rd_skid2_2_vld;
  assign _2159_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) _1285_;
  assign _2160_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) rd_take_n_dly[2];
  assign _2161_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) cq_rd_credit[2];
  assign _2162_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) cq_rd2_prdy_d;
  assign _2163_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) _1305_;
  assign _2164_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) rd_skid3_0_vld;
  assign _2165_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) rd_skid3_1_vld;
  assign _2166_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *) rd_skid3_2_vld;
  assign _2167_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) _1308_;
  assign _2168_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) rd_take_n_dly[3];
  assign _2169_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) cq_rd_credit[3];
  assign _2170_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) cq_rd3_prdy_d;
  assign _2171_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) _1329_;
  assign _2172_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) rd_skid4_0_vld;
  assign _2173_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) rd_skid4_1_vld;
  assign _2174_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *) rd_skid4_2_vld;
  assign _2175_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) _1332_;
  assign _2176_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) rd_take_n_dly[4];
  assign _2177_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) cq_rd_credit[4];
  assign _2178_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) cq_rd4_prdy_d;
  assign _2179_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) _1353_;
  assign _2180_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) rd_skid5_0_vld;
  assign _2181_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) rd_skid5_1_vld;
  assign _2182_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *) rd_skid5_2_vld;
  assign _2183_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) _1356_;
  assign _2184_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) rd_take_n_dly[5];
  assign _2185_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) cq_rd_credit[5];
  assign _2186_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) cq_rd5_prdy_d;
  assign _2187_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) _1376_;
  assign _2188_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) rd_skid6_0_vld;
  assign _2189_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) rd_skid6_1_vld;
  assign _2190_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *) rd_skid6_2_vld;
  assign _2191_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) _1380_;
  assign _2192_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) rd_take_n_dly[6];
  assign _2193_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) cq_rd_credit[6];
  assign _2194_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) cq_rd6_prdy_d;
  assign _2195_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) _1400_;
  assign _2196_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) rd_skid7_0_vld;
  assign _2197_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) rd_skid7_1_vld;
  assign _2198_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *) rd_skid7_2_vld;
  assign _2199_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) _1404_;
  assign _2200_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) rd_take_n_dly[7];
  assign _2201_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) cq_rd_credit[7];
  assign _2202_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) cq_rd7_prdy_d;
  assign _2203_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) _1424_;
  assign _2204_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) rd_skid8_0_vld;
  assign _2205_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) rd_skid8_1_vld;
  assign _2206_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *) rd_skid8_2_vld;
  assign _2207_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) _1427_;
  assign _2208_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) rd_take_n_dly[8];
  assign _2209_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) cq_rd_credit[8];
  assign _2210_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) cq_rd8_prdy_d;
  assign _2211_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) _1448_;
  assign _2212_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) rd_skid9_0_vld;
  assign _2213_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) rd_skid9_1_vld;
  assign _2214_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *) rd_skid9_2_vld;
  assign _2215_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) _1451_;
  assign _2216_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) rd_take_n_dly[9];
  assign _2217_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) cq_rd_credit[9];
  assign _2218_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) cq_rd9_prdy_d;
  assign _2219_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) _1472_;
  assign _2220_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3513" *) cq_rd_take_elig[0];
  assign _2221_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3514" *) cq_rd_take_elig[9];
  assign _2222_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3515" *) cq_rd_take_elig[8];
  assign _2223_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3516" *) cq_rd_take_elig[7];
  assign _2224_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3517" *) cq_rd_take_elig[6];
  assign _2225_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3518" *) cq_rd_take_elig[5];
  assign _2226_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3519" *) cq_rd_take_elig[4];
  assign _2227_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3520" *) cq_rd_take_elig[3];
  assign _2228_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3521" *) cq_rd_take_elig[2];
  assign _2229_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3524" *) cq_rd_take_elig[1];
  assign _2230_ = rd_pushing || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing_q;
  assign update_rd_take_n_dly = cq_rd_take || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2069" *) rd_take_dly;
  assign _2231_ = rd_take_dly || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:211" *) rd_pushing;
  assign _2232_ = rd_pushing || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2264" *) cq_rd_take;
  assign _2233_ = _1165_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *) _1167_;
  assign _2234_ = _1169_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *) _1171_;
  assign _2235_ = _1173_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *) _1175_;
  assign _2236_ = _1176_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *) _1178_;
  assign _2237_ = _1180_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *) _1182_;
  assign _2238_ = _1184_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *) _1186_;
  assign _2239_ = _1187_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *) _1189_;
  assign _2240_ = _1191_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *) _1193_;
  assign _2241_ = _1194_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *) _1196_;
  assign _2242_ = _1198_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *) _1200_;
  assign cq_rd0_pvld = rd_skid0_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2566" *) rd_pre_bypassing0;
  assign _2243_ = rd_bypassing0 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) rd_take_n_dly[0];
  assign _2244_ = _2140_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) _1238_;
  assign _2245_ = _2141_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *) _1241_;
  assign _2246_ = rd_skid0_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) _2143_;
  assign _2247_ = rd_skid0_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) _1248_;
  assign _2248_ = _2247_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) rd_take_n_dly[0];
  assign _2249_ = rd_skid0_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) rd_bypassing0;
  assign _2250_ = _2249_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) rd_take_n_dly[0];
  assign _2251_ = rd_skid0_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *) _1250_;
  assign _2252_ = rd_skid0_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *) _1245_;
  assign _2253_ = cq_rd0_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) _2140_;
  assign _2254_ = _2253_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) _2141_;
  assign _2255_ = _2254_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) _1252_;
  assign _2256_ = cq_rd_credit[0] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2624" *) cq_rd0_credits_ne0;
  assign _2257_ = _2144_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2626" *) rd_skid0_0_vld;
  assign _2258_ = _2142_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) _2141_;
  assign _2259_ = _2258_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2627" *) _2147_;
  assign cq_rd1_pvld = rd_skid1_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2662" *) rd_pre_bypassing1;
  assign _2260_ = rd_bypassing1 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) rd_take_n_dly[1];
  assign _2261_ = _2148_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) _1262_;
  assign _2262_ = _2149_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *) _1265_;
  assign _2263_ = rd_skid1_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) _2151_;
  assign _2264_ = rd_skid1_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) _1272_;
  assign _2265_ = _2264_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) rd_take_n_dly[1];
  assign _2266_ = rd_skid1_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) rd_bypassing1;
  assign _2267_ = _2266_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) rd_take_n_dly[1];
  assign _2268_ = rd_skid1_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *) _1273_;
  assign _2269_ = rd_skid1_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *) _1268_;
  assign _2270_ = cq_rd1_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) _2148_;
  assign _2271_ = _2270_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) _2149_;
  assign _2272_ = _2271_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) _1276_;
  assign _2273_ = cq_rd_credit[1] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2720" *) cq_rd1_credits_ne0;
  assign _2274_ = _2152_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2722" *) rd_skid1_0_vld;
  assign _2275_ = _2150_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) _2149_;
  assign _2276_ = _2275_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2723" *) _2155_;
  assign cq_rd2_pvld = rd_skid2_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2758" *) rd_pre_bypassing2;
  assign _2277_ = rd_bypassing2 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) rd_take_n_dly[2];
  assign _2278_ = _2156_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) _1286_;
  assign _2279_ = _2157_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *) _1289_;
  assign _2280_ = rd_skid2_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) _2159_;
  assign _2281_ = rd_skid2_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) _1296_;
  assign _2282_ = _2281_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) rd_take_n_dly[2];
  assign _2283_ = rd_skid2_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) rd_bypassing2;
  assign _2284_ = _2283_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) rd_take_n_dly[2];
  assign _2285_ = rd_skid2_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *) _1297_;
  assign _2286_ = rd_skid2_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *) _1292_;
  assign _2287_ = cq_rd2_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) _2156_;
  assign _2288_ = _2287_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) _2157_;
  assign _2289_ = _2288_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) _1300_;
  assign _2290_ = cq_rd_credit[2] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2816" *) cq_rd2_credits_ne0;
  assign _2291_ = _2160_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2818" *) rd_skid2_0_vld;
  assign _2292_ = _2158_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) _2157_;
  assign _2293_ = _2292_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2819" *) _2163_;
  assign cq_rd3_pvld = rd_skid3_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2854" *) rd_pre_bypassing3;
  assign _2294_ = rd_bypassing3 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) rd_take_n_dly[3];
  assign _2295_ = _2164_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) _1309_;
  assign _2296_ = _2165_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *) _1313_;
  assign _2297_ = rd_skid3_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) _2167_;
  assign _2298_ = rd_skid3_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) _1320_;
  assign _2299_ = _2298_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) rd_take_n_dly[3];
  assign _2300_ = rd_skid3_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) rd_bypassing3;
  assign _2301_ = _2300_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) rd_take_n_dly[3];
  assign _2302_ = rd_skid3_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *) _1321_;
  assign _2303_ = rd_skid3_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *) _1316_;
  assign _2304_ = cq_rd3_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) _2164_;
  assign _2305_ = _2304_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) _2165_;
  assign _2306_ = _2305_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) _1324_;
  assign _2307_ = cq_rd_credit[3] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2912" *) cq_rd3_credits_ne0;
  assign _2308_ = _2168_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2914" *) rd_skid3_0_vld;
  assign _2309_ = _2166_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) _2165_;
  assign _2310_ = _2309_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2915" *) _2171_;
  assign cq_rd4_pvld = rd_skid4_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2950" *) rd_pre_bypassing4;
  assign _2311_ = rd_bypassing4 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) rd_take_n_dly[4];
  assign _2312_ = _2172_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) _1333_;
  assign _2313_ = _2173_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *) _1337_;
  assign _2314_ = rd_skid4_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) _2175_;
  assign _2315_ = rd_skid4_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) _1344_;
  assign _2316_ = _2315_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) rd_take_n_dly[4];
  assign _2317_ = rd_skid4_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) rd_bypassing4;
  assign _2318_ = _2317_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) rd_take_n_dly[4];
  assign _2319_ = rd_skid4_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *) _1345_;
  assign _2320_ = rd_skid4_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *) _1340_;
  assign _2321_ = cq_rd4_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) _2172_;
  assign _2322_ = _2321_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) _2173_;
  assign _2323_ = _2322_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) _1347_;
  assign _2324_ = cq_rd_credit[4] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3008" *) cq_rd4_credits_ne0;
  assign _2325_ = _2176_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3010" *) rd_skid4_0_vld;
  assign _2326_ = _2174_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) _2173_;
  assign _2327_ = _2326_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3011" *) _2179_;
  assign cq_rd5_pvld = rd_skid5_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3046" *) rd_pre_bypassing5;
  assign _2328_ = rd_bypassing5 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) rd_take_n_dly[5];
  assign _2329_ = _2180_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) _1357_;
  assign _2330_ = _2181_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *) _1361_;
  assign _2331_ = rd_skid5_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) _2183_;
  assign _2332_ = rd_skid5_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) _1367_;
  assign _2333_ = _2332_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) rd_take_n_dly[5];
  assign _2334_ = rd_skid5_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) rd_bypassing5;
  assign _2335_ = _2334_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) rd_take_n_dly[5];
  assign _2336_ = rd_skid5_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *) _1369_;
  assign _2337_ = rd_skid5_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *) _1364_;
  assign _2338_ = cq_rd5_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) _2180_;
  assign _2339_ = _2338_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) _2181_;
  assign _2340_ = _2339_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) _1371_;
  assign _2341_ = cq_rd_credit[5] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3104" *) cq_rd5_credits_ne0;
  assign _2342_ = _2184_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3106" *) rd_skid5_0_vld;
  assign _2343_ = _2182_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) _2181_;
  assign _2344_ = _2343_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3107" *) _2187_;
  assign cq_rd6_pvld = rd_skid6_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3142" *) rd_pre_bypassing6;
  assign _2345_ = rd_bypassing6 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) rd_take_n_dly[6];
  assign _2346_ = _2188_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) _1381_;
  assign _2347_ = _2189_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *) _1384_;
  assign _2348_ = rd_skid6_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) _2191_;
  assign _2349_ = rd_skid6_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) _1391_;
  assign _2350_ = _2349_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) rd_take_n_dly[6];
  assign _2351_ = rd_skid6_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) rd_bypassing6;
  assign _2352_ = _2351_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) rd_take_n_dly[6];
  assign _2353_ = rd_skid6_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *) _1392_;
  assign _2354_ = rd_skid6_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *) _1388_;
  assign _2355_ = cq_rd6_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) _2188_;
  assign _2356_ = _2355_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) _2189_;
  assign _2357_ = _2356_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) _1395_;
  assign _2358_ = cq_rd_credit[6] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3200" *) cq_rd6_credits_ne0;
  assign _2359_ = _2192_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3202" *) rd_skid6_0_vld;
  assign _2360_ = _2190_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) _2189_;
  assign _2361_ = _2360_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3203" *) _2195_;
  assign cq_rd7_pvld = rd_skid7_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3238" *) rd_pre_bypassing7;
  assign _2362_ = rd_bypassing7 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) rd_take_n_dly[7];
  assign _2363_ = _2196_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) _1405_;
  assign _2364_ = _2197_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *) _1408_;
  assign _2365_ = rd_skid7_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) _2199_;
  assign _2366_ = rd_skid7_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) _1415_;
  assign _2367_ = _2366_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) rd_take_n_dly[7];
  assign _2368_ = rd_skid7_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) rd_bypassing7;
  assign _2369_ = _2368_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) rd_take_n_dly[7];
  assign _2370_ = rd_skid7_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *) _1416_;
  assign _2371_ = rd_skid7_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *) _1412_;
  assign _2372_ = cq_rd7_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) _2196_;
  assign _2373_ = _2372_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) _2197_;
  assign _2374_ = _2373_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) _1419_;
  assign _2375_ = cq_rd_credit[7] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3296" *) cq_rd7_credits_ne0;
  assign _2376_ = _2200_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3298" *) rd_skid7_0_vld;
  assign _2377_ = _2198_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) _2197_;
  assign _2378_ = _2377_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3299" *) _2203_;
  assign cq_rd8_pvld = rd_skid8_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3334" *) rd_pre_bypassing8;
  assign _2379_ = rd_bypassing8 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) rd_take_n_dly[8];
  assign _2380_ = _2204_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) _1428_;
  assign _2381_ = _2205_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *) _1432_;
  assign _2382_ = rd_skid8_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) _2207_;
  assign _2383_ = rd_skid8_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) _1439_;
  assign _2384_ = _2383_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) rd_take_n_dly[8];
  assign _2385_ = rd_skid8_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) rd_bypassing8;
  assign _2386_ = _2385_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) rd_take_n_dly[8];
  assign _2387_ = rd_skid8_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *) _1440_;
  assign _2388_ = rd_skid8_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *) _1436_;
  assign _2389_ = cq_rd8_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) _2204_;
  assign _2390_ = _2389_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) _2205_;
  assign _2391_ = _2390_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) _1443_;
  assign _2392_ = cq_rd_credit[8] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3392" *) cq_rd8_credits_ne0;
  assign _2393_ = _2208_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3394" *) rd_skid8_0_vld;
  assign _2394_ = _2206_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) _2205_;
  assign _2395_ = _2394_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3395" *) _2211_;
  assign cq_rd9_pvld = rd_skid9_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3430" *) rd_pre_bypassing9;
  assign _2396_ = rd_bypassing9 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) rd_take_n_dly[9];
  assign _2397_ = _2212_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) _1452_;
  assign _2398_ = _2213_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *) _1456_;
  assign _2399_ = rd_skid9_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) _2215_;
  assign _2400_ = rd_skid9_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) _1463_;
  assign _2401_ = _2400_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) rd_take_n_dly[9];
  assign _2402_ = rd_skid9_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) rd_bypassing9;
  assign _2403_ = _2402_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) rd_take_n_dly[9];
  assign _2404_ = rd_skid9_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *) _1464_;
  assign _2405_ = rd_skid9_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *) _1459_;
  assign _2406_ = cq_rd9_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) _2212_;
  assign _2407_ = _2406_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) _2213_;
  assign _2408_ = _2407_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) _1466_;
  assign _2409_ = cq_rd_credit[9] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3488" *) cq_rd9_credits_ne0;
  assign _2410_ = _2216_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3490" *) rd_skid9_0_vld;
  assign _2411_ = _2214_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) _2213_;
  assign _2412_ = _2411_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3491" *) _2219_;
  assign _2413_ = rd_bypassing0 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing1;
  assign _2414_ = _2413_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing2;
  assign _2415_ = _2414_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing3;
  assign _2416_ = _2415_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing4;
  assign _2417_ = _2416_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing5;
  assign _2418_ = _2417_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing6;
  assign _2419_ = _2418_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing7;
  assign _2420_ = _2419_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing8;
  assign wr_bypassing = _2420_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3630" *) rd_bypassing9;
  assign _2421_ = wr_reserving || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) rd_pushing;
  assign _2422_ = _2421_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) rd_take_dly;
  assign _2423_ = _2422_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) wr_reserving;
  assign _2424_ = _2423_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) _2477_;
  assign _2425_ = _2424_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) rd_take_dly;
  assign _2426_ = _2232_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) _2478_;
  assign _2427_ = _2426_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) rd_take_dly;
  assign nvdla_core_clk_mgated_enable = _2425_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) _2427_;
  assign _2428_ = nvdla_core_clk_mgated_enable || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1237_;
  assign _2429_ = _2428_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing0;
  assign _2430_ = _2429_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1261_;
  assign _2431_ = _2430_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing1;
  assign _2432_ = _2431_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1285_;
  assign _2433_ = _2432_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing2;
  assign _2434_ = _2433_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1308_;
  assign _2435_ = _2434_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing3;
  assign _2436_ = _2435_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1332_;
  assign _2437_ = _2436_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing4;
  assign _2438_ = _2437_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1356_;
  assign _2439_ = _2438_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing5;
  assign _2440_ = _2439_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1380_;
  assign _2441_ = _2440_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing6;
  assign _2442_ = _2441_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1404_;
  assign _2443_ = _2442_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing7;
  assign _2444_ = _2443_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1427_;
  assign _2445_ = _2444_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) rd_bypassing8;
  assign _2446_ = _2445_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3665" *) _1451_;
  assign nvdla_core_clk_mgated_skid_enable = _2446_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3676" *) rd_bypassing9;
  assign _2447_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2457" *) cq_rd_count0;
  assign _2448_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2458" *) cq_rd_count1;
  assign _2449_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2459" *) cq_rd_count2;
  assign _2450_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2460" *) cq_rd_count3;
  assign _2451_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2461" *) cq_rd_count4;
  assign _2452_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2462" *) cq_rd_count5;
  assign _2453_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2463" *) cq_rd_count6;
  assign _2454_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2464" *) cq_rd_count7;
  assign _2455_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2465" *) cq_rd_count8;
  assign _2456_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2466" *) cq_rd_count9;
  assign _2457_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *) cq_rd0_credits_w_take_next;
  assign _2458_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *) cq_rd0_credits_wo_take_next;
  assign _2459_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *) cq_rd1_credits_w_take_next;
  assign _2460_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *) cq_rd1_credits_wo_take_next;
  assign _2461_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *) cq_rd2_credits_w_take_next;
  assign _2462_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *) cq_rd2_credits_wo_take_next;
  assign _2463_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *) cq_rd3_credits_w_take_next;
  assign _2464_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *) cq_rd3_credits_wo_take_next;
  assign _2465_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *) cq_rd4_credits_w_take_next;
  assign _2466_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *) cq_rd4_credits_wo_take_next;
  assign _2467_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *) cq_rd5_credits_w_take_next;
  assign _2468_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *) cq_rd5_credits_wo_take_next;
  assign _2469_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *) cq_rd6_credits_w_take_next;
  assign _2470_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *) cq_rd6_credits_wo_take_next;
  assign _2471_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *) cq_rd7_credits_w_take_next;
  assign _2472_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *) cq_rd7_credits_wo_take_next;
  assign _2473_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *) cq_rd8_credits_w_take_next;
  assign _2474_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *) cq_rd8_credits_wo_take_next;
  assign _2475_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *) cq_rd9_credits_w_take_next;
  assign _2476_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *) cq_rd9_credits_wo_take_next;
  assign _2477_ = cq_wr_busy_int != (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) cq_wr_busy_next;
  assign _2478_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3653" *) cq_rd_credit;
  assign flag_l0_0 = free_adr_mask[1] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1500" *) free_adr_mask[0];
  assign flag_l0_1 = free_adr_mask[3] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1501" *) free_adr_mask[2];
  assign flag_l0_2 = free_adr_mask[5] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1502" *) free_adr_mask[4];
  assign flag_l0_3 = free_adr_mask[7] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1503" *) free_adr_mask[6];
  assign flag_l0_4 = free_adr_mask[9] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1504" *) free_adr_mask[8];
  assign flag_l0_5 = free_adr_mask[11] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1505" *) free_adr_mask[10];
  assign flag_l0_6 = free_adr_mask[13] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1506" *) free_adr_mask[12];
  assign flag_l0_7 = free_adr_mask[15] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1507" *) free_adr_mask[14];
  assign flag_l0_8 = free_adr_mask[17] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1508" *) free_adr_mask[16];
  assign flag_l0_9 = free_adr_mask[19] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1509" *) free_adr_mask[18];
  assign flag_l0_10 = free_adr_mask[21] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1510" *) free_adr_mask[20];
  assign flag_l0_11 = free_adr_mask[23] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1511" *) free_adr_mask[22];
  assign flag_l0_12 = free_adr_mask[25] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1512" *) free_adr_mask[24];
  assign flag_l0_13 = free_adr_mask[27] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1513" *) free_adr_mask[26];
  assign flag_l0_14 = free_adr_mask[29] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1514" *) free_adr_mask[28];
  assign flag_l0_15 = free_adr_mask[31] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1515" *) free_adr_mask[30];
  assign flag_l0_16 = free_adr_mask[33] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1516" *) free_adr_mask[32];
  assign flag_l0_17 = free_adr_mask[35] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1517" *) free_adr_mask[34];
  assign flag_l0_18 = free_adr_mask[37] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1518" *) free_adr_mask[36];
  assign flag_l0_19 = free_adr_mask[39] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1519" *) free_adr_mask[38];
  assign flag_l0_20 = free_adr_mask[41] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1520" *) free_adr_mask[40];
  assign flag_l0_21 = free_adr_mask[43] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1521" *) free_adr_mask[42];
  assign flag_l0_22 = free_adr_mask[45] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1522" *) free_adr_mask[44];
  assign flag_l0_23 = free_adr_mask[47] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1523" *) free_adr_mask[46];
  assign flag_l0_24 = free_adr_mask[49] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1524" *) free_adr_mask[48];
  assign flag_l0_25 = free_adr_mask[51] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1525" *) free_adr_mask[50];
  assign flag_l0_26 = free_adr_mask[53] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1526" *) free_adr_mask[52];
  assign flag_l0_27 = free_adr_mask[55] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1527" *) free_adr_mask[54];
  assign flag_l0_28 = free_adr_mask[57] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1528" *) free_adr_mask[56];
  assign flag_l0_29 = free_adr_mask[59] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1529" *) free_adr_mask[58];
  assign flag_l0_30 = free_adr_mask[61] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1530" *) free_adr_mask[60];
  assign flag_l0_31 = free_adr_mask[63] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1531" *) free_adr_mask[62];
  assign flag_l0_32 = free_adr_mask[65] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1532" *) free_adr_mask[64];
  assign flag_l0_33 = free_adr_mask[67] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1533" *) free_adr_mask[66];
  assign flag_l0_34 = free_adr_mask[69] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1534" *) free_adr_mask[68];
  assign flag_l0_35 = free_adr_mask[71] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1535" *) free_adr_mask[70];
  assign flag_l0_36 = free_adr_mask[73] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1536" *) free_adr_mask[72];
  assign flag_l0_37 = free_adr_mask[75] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1537" *) free_adr_mask[74];
  assign flag_l0_38 = free_adr_mask[77] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1538" *) free_adr_mask[76];
  assign flag_l0_39 = free_adr_mask[79] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1539" *) free_adr_mask[78];
  assign flag_l0_40 = free_adr_mask[81] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1540" *) free_adr_mask[80];
  assign flag_l0_41 = free_adr_mask[83] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1541" *) free_adr_mask[82];
  assign flag_l0_42 = free_adr_mask[85] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1542" *) free_adr_mask[84];
  assign flag_l0_43 = free_adr_mask[87] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1543" *) free_adr_mask[86];
  assign flag_l0_44 = free_adr_mask[89] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1544" *) free_adr_mask[88];
  assign flag_l0_45 = free_adr_mask[91] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1545" *) free_adr_mask[90];
  assign flag_l0_46 = free_adr_mask[93] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1546" *) free_adr_mask[92];
  assign flag_l0_47 = free_adr_mask[95] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1547" *) free_adr_mask[94];
  assign flag_l0_48 = free_adr_mask[97] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1548" *) free_adr_mask[96];
  assign flag_l0_49 = free_adr_mask[99] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1549" *) free_adr_mask[98];
  assign flag_l0_50 = free_adr_mask[101] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1550" *) free_adr_mask[100];
  assign flag_l0_51 = free_adr_mask[103] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1551" *) free_adr_mask[102];
  assign flag_l0_52 = free_adr_mask[105] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1552" *) free_adr_mask[104];
  assign flag_l0_53 = free_adr_mask[107] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1553" *) free_adr_mask[106];
  assign flag_l0_54 = free_adr_mask[109] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1554" *) free_adr_mask[108];
  assign flag_l0_55 = free_adr_mask[111] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1555" *) free_adr_mask[110];
  assign flag_l0_56 = free_adr_mask[113] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1556" *) free_adr_mask[112];
  assign flag_l0_57 = free_adr_mask[115] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1557" *) free_adr_mask[114];
  assign flag_l0_58 = free_adr_mask[117] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1558" *) free_adr_mask[116];
  assign flag_l0_59 = free_adr_mask[119] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1559" *) free_adr_mask[118];
  assign flag_l0_60 = free_adr_mask[121] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1560" *) free_adr_mask[120];
  assign flag_l0_61 = free_adr_mask[123] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1561" *) free_adr_mask[122];
  assign flag_l0_62 = free_adr_mask[125] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1562" *) free_adr_mask[124];
  assign flag_l0_63 = free_adr_mask[127] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1563" *) free_adr_mask[126];
  assign flag_l0_64 = free_adr_mask[129] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1564" *) free_adr_mask[128];
  assign flag_l0_65 = free_adr_mask[131] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1565" *) free_adr_mask[130];
  assign flag_l0_66 = free_adr_mask[133] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1566" *) free_adr_mask[132];
  assign flag_l0_67 = free_adr_mask[135] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1567" *) free_adr_mask[134];
  assign flag_l0_68 = free_adr_mask[137] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1568" *) free_adr_mask[136];
  assign flag_l0_69 = free_adr_mask[139] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1569" *) free_adr_mask[138];
  assign flag_l0_70 = free_adr_mask[141] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1570" *) free_adr_mask[140];
  assign flag_l0_71 = free_adr_mask[143] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1571" *) free_adr_mask[142];
  assign flag_l0_72 = free_adr_mask[145] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1572" *) free_adr_mask[144];
  assign flag_l0_73 = free_adr_mask[147] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1573" *) free_adr_mask[146];
  assign flag_l0_74 = free_adr_mask[149] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1574" *) free_adr_mask[148];
  assign flag_l0_75 = free_adr_mask[151] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1575" *) free_adr_mask[150];
  assign flag_l0_76 = free_adr_mask[153] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1576" *) free_adr_mask[152];
  assign flag_l0_77 = free_adr_mask[155] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1577" *) free_adr_mask[154];
  assign flag_l0_78 = free_adr_mask[157] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1578" *) free_adr_mask[156];
  assign flag_l0_79 = free_adr_mask[159] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1579" *) free_adr_mask[158];
  assign flag_l0_80 = free_adr_mask[161] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1580" *) free_adr_mask[160];
  assign flag_l0_81 = free_adr_mask[163] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1581" *) free_adr_mask[162];
  assign flag_l0_82 = free_adr_mask[165] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1582" *) free_adr_mask[164];
  assign flag_l0_83 = free_adr_mask[167] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1583" *) free_adr_mask[166];
  assign flag_l0_84 = free_adr_mask[169] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1584" *) free_adr_mask[168];
  assign flag_l0_85 = free_adr_mask[171] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1585" *) free_adr_mask[170];
  assign flag_l0_86 = free_adr_mask[173] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1586" *) free_adr_mask[172];
  assign flag_l0_87 = free_adr_mask[175] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1587" *) free_adr_mask[174];
  assign flag_l0_88 = free_adr_mask[177] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1588" *) free_adr_mask[176];
  assign flag_l0_89 = free_adr_mask[179] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1589" *) free_adr_mask[178];
  assign flag_l0_90 = free_adr_mask[181] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1590" *) free_adr_mask[180];
  assign flag_l0_91 = free_adr_mask[183] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1591" *) free_adr_mask[182];
  assign flag_l0_92 = free_adr_mask[185] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1592" *) free_adr_mask[184];
  assign flag_l0_93 = free_adr_mask[187] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1593" *) free_adr_mask[186];
  assign flag_l0_94 = free_adr_mask[189] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1594" *) free_adr_mask[188];
  assign flag_l0_95 = free_adr_mask[191] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1595" *) free_adr_mask[190];
  assign flag_l0_96 = free_adr_mask[193] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1596" *) free_adr_mask[192];
  assign flag_l0_97 = free_adr_mask[195] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1597" *) free_adr_mask[194];
  assign flag_l0_98 = free_adr_mask[197] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1598" *) free_adr_mask[196];
  assign flag_l0_99 = free_adr_mask[199] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1599" *) free_adr_mask[198];
  assign flag_l0_100 = free_adr_mask[201] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1600" *) free_adr_mask[200];
  assign flag_l0_101 = free_adr_mask[203] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1601" *) free_adr_mask[202];
  assign flag_l0_102 = free_adr_mask[205] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1602" *) free_adr_mask[204];
  assign flag_l0_103 = free_adr_mask[207] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1603" *) free_adr_mask[206];
  assign flag_l0_104 = free_adr_mask[209] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1604" *) free_adr_mask[208];
  assign flag_l0_105 = free_adr_mask[211] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1605" *) free_adr_mask[210];
  assign flag_l0_106 = free_adr_mask[213] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1606" *) free_adr_mask[212];
  assign flag_l0_107 = free_adr_mask[215] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1607" *) free_adr_mask[214];
  assign flag_l0_108 = free_adr_mask[217] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1608" *) free_adr_mask[216];
  assign flag_l0_109 = free_adr_mask[219] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1609" *) free_adr_mask[218];
  assign flag_l0_110 = free_adr_mask[221] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1610" *) free_adr_mask[220];
  assign flag_l0_111 = free_adr_mask[223] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1611" *) free_adr_mask[222];
  assign flag_l0_112 = free_adr_mask[225] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1612" *) free_adr_mask[224];
  assign flag_l0_113 = free_adr_mask[227] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1613" *) free_adr_mask[226];
  assign flag_l0_114 = free_adr_mask[229] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1614" *) free_adr_mask[228];
  assign flag_l0_115 = free_adr_mask[231] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1615" *) free_adr_mask[230];
  assign flag_l0_116 = free_adr_mask[233] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1616" *) free_adr_mask[232];
  assign flag_l0_117 = free_adr_mask[235] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1617" *) free_adr_mask[234];
  assign flag_l0_118 = free_adr_mask[237] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1618" *) free_adr_mask[236];
  assign flag_l0_119 = free_adr_mask[239] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1619" *) free_adr_mask[238];
  assign flag_l0_120 = free_adr_mask[241] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1620" *) free_adr_mask[240];
  assign flag_l0_121 = free_adr_mask[243] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1621" *) free_adr_mask[242];
  assign flag_l0_122 = free_adr_mask[245] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1622" *) free_adr_mask[244];
  assign flag_l0_123 = free_adr_mask[247] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1623" *) free_adr_mask[246];
  assign flag_l0_124 = free_adr_mask[249] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1624" *) free_adr_mask[248];
  assign flag_l0_125 = free_adr_mask[251] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1625" *) free_adr_mask[250];
  assign flag_l0_126 = free_adr_mask[253] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1626" *) free_adr_mask[252];
  assign flag_l1_0 = flag_l0_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1627" *) flag_l0_0;
  assign flag_l1_1 = flag_l0_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1628" *) flag_l0_2;
  assign flag_l1_2 = flag_l0_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1629" *) flag_l0_4;
  assign flag_l1_3 = flag_l0_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1630" *) flag_l0_6;
  assign flag_l1_4 = flag_l0_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1631" *) flag_l0_8;
  assign flag_l1_5 = flag_l0_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1632" *) flag_l0_10;
  assign flag_l1_6 = flag_l0_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1633" *) flag_l0_12;
  assign flag_l1_7 = flag_l0_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1634" *) flag_l0_14;
  assign flag_l1_8 = flag_l0_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1635" *) flag_l0_16;
  assign flag_l1_9 = flag_l0_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1636" *) flag_l0_18;
  assign flag_l1_10 = flag_l0_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1637" *) flag_l0_20;
  assign flag_l1_11 = flag_l0_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1638" *) flag_l0_22;
  assign flag_l1_12 = flag_l0_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1639" *) flag_l0_24;
  assign flag_l1_13 = flag_l0_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1640" *) flag_l0_26;
  assign flag_l1_14 = flag_l0_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1641" *) flag_l0_28;
  assign flag_l1_15 = flag_l0_31 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1642" *) flag_l0_30;
  assign flag_l1_16 = flag_l0_33 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1643" *) flag_l0_32;
  assign flag_l1_17 = flag_l0_35 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1644" *) flag_l0_34;
  assign flag_l1_18 = flag_l0_37 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1645" *) flag_l0_36;
  assign flag_l1_19 = flag_l0_39 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1646" *) flag_l0_38;
  assign flag_l1_20 = flag_l0_41 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1647" *) flag_l0_40;
  assign flag_l1_21 = flag_l0_43 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1648" *) flag_l0_42;
  assign flag_l1_22 = flag_l0_45 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1649" *) flag_l0_44;
  assign flag_l1_23 = flag_l0_47 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1650" *) flag_l0_46;
  assign flag_l1_24 = flag_l0_49 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1651" *) flag_l0_48;
  assign flag_l1_25 = flag_l0_51 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1652" *) flag_l0_50;
  assign flag_l1_26 = flag_l0_53 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1653" *) flag_l0_52;
  assign flag_l1_27 = flag_l0_55 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1654" *) flag_l0_54;
  assign flag_l1_28 = flag_l0_57 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1655" *) flag_l0_56;
  assign flag_l1_29 = flag_l0_59 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1656" *) flag_l0_58;
  assign flag_l1_30 = flag_l0_61 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1657" *) flag_l0_60;
  assign flag_l1_31 = flag_l0_63 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1658" *) flag_l0_62;
  assign flag_l1_32 = flag_l0_65 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1659" *) flag_l0_64;
  assign flag_l1_33 = flag_l0_67 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1660" *) flag_l0_66;
  assign flag_l1_34 = flag_l0_69 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1661" *) flag_l0_68;
  assign flag_l1_35 = flag_l0_71 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1662" *) flag_l0_70;
  assign flag_l1_36 = flag_l0_73 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1663" *) flag_l0_72;
  assign flag_l1_37 = flag_l0_75 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1664" *) flag_l0_74;
  assign flag_l1_38 = flag_l0_77 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1665" *) flag_l0_76;
  assign flag_l1_39 = flag_l0_79 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1666" *) flag_l0_78;
  assign flag_l1_40 = flag_l0_81 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1667" *) flag_l0_80;
  assign flag_l1_41 = flag_l0_83 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1668" *) flag_l0_82;
  assign flag_l1_42 = flag_l0_85 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1669" *) flag_l0_84;
  assign flag_l1_43 = flag_l0_87 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1670" *) flag_l0_86;
  assign flag_l1_44 = flag_l0_89 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1671" *) flag_l0_88;
  assign flag_l1_45 = flag_l0_91 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1672" *) flag_l0_90;
  assign flag_l1_46 = flag_l0_93 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1673" *) flag_l0_92;
  assign flag_l1_47 = flag_l0_95 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1674" *) flag_l0_94;
  assign flag_l1_48 = flag_l0_97 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1675" *) flag_l0_96;
  assign flag_l1_49 = flag_l0_99 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1676" *) flag_l0_98;
  assign flag_l1_50 = flag_l0_101 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1677" *) flag_l0_100;
  assign flag_l1_51 = flag_l0_103 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1678" *) flag_l0_102;
  assign flag_l1_52 = flag_l0_105 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1679" *) flag_l0_104;
  assign flag_l1_53 = flag_l0_107 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1680" *) flag_l0_106;
  assign flag_l1_54 = flag_l0_109 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1681" *) flag_l0_108;
  assign flag_l1_55 = flag_l0_111 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1682" *) flag_l0_110;
  assign flag_l1_56 = flag_l0_113 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1683" *) flag_l0_112;
  assign flag_l1_57 = flag_l0_115 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1684" *) flag_l0_114;
  assign flag_l1_58 = flag_l0_117 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1685" *) flag_l0_116;
  assign flag_l1_59 = flag_l0_119 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1686" *) flag_l0_118;
  assign flag_l1_60 = flag_l0_121 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1687" *) flag_l0_120;
  assign flag_l1_61 = flag_l0_123 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1688" *) flag_l0_122;
  assign flag_l1_62 = flag_l0_125 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1689" *) flag_l0_124;
  assign flag_l2_0 = flag_l1_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1690" *) flag_l1_0;
  assign flag_l2_1 = flag_l1_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1691" *) flag_l1_2;
  assign flag_l2_2 = flag_l1_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1692" *) flag_l1_4;
  assign flag_l2_3 = flag_l1_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1693" *) flag_l1_6;
  assign flag_l2_4 = flag_l1_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1694" *) flag_l1_8;
  assign flag_l2_5 = flag_l1_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1695" *) flag_l1_10;
  assign flag_l2_6 = flag_l1_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1696" *) flag_l1_12;
  assign flag_l2_7 = flag_l1_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1697" *) flag_l1_14;
  assign flag_l2_8 = flag_l1_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1698" *) flag_l1_16;
  assign flag_l2_9 = flag_l1_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1699" *) flag_l1_18;
  assign flag_l2_10 = flag_l1_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1700" *) flag_l1_20;
  assign flag_l2_11 = flag_l1_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1701" *) flag_l1_22;
  assign flag_l2_12 = flag_l1_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1702" *) flag_l1_24;
  assign flag_l2_13 = flag_l1_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1703" *) flag_l1_26;
  assign flag_l2_14 = flag_l1_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1704" *) flag_l1_28;
  assign flag_l2_15 = flag_l1_31 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1705" *) flag_l1_30;
  assign flag_l2_16 = flag_l1_33 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1706" *) flag_l1_32;
  assign flag_l2_17 = flag_l1_35 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1707" *) flag_l1_34;
  assign flag_l2_18 = flag_l1_37 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1708" *) flag_l1_36;
  assign flag_l2_19 = flag_l1_39 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1709" *) flag_l1_38;
  assign flag_l2_20 = flag_l1_41 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1710" *) flag_l1_40;
  assign flag_l2_21 = flag_l1_43 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1711" *) flag_l1_42;
  assign flag_l2_22 = flag_l1_45 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1712" *) flag_l1_44;
  assign flag_l2_23 = flag_l1_47 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1713" *) flag_l1_46;
  assign flag_l2_24 = flag_l1_49 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1714" *) flag_l1_48;
  assign flag_l2_25 = flag_l1_51 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1715" *) flag_l1_50;
  assign flag_l2_26 = flag_l1_53 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1716" *) flag_l1_52;
  assign flag_l2_27 = flag_l1_55 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1717" *) flag_l1_54;
  assign flag_l2_28 = flag_l1_57 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1718" *) flag_l1_56;
  assign flag_l2_29 = flag_l1_59 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1719" *) flag_l1_58;
  assign flag_l2_30 = flag_l1_61 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1720" *) flag_l1_60;
  assign flag_l3_0 = flag_l2_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1721" *) flag_l2_0;
  assign flag_l3_1 = flag_l2_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1722" *) flag_l2_2;
  assign flag_l3_2 = flag_l2_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1723" *) flag_l2_4;
  assign flag_l3_3 = flag_l2_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1724" *) flag_l2_6;
  assign flag_l3_4 = flag_l2_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1725" *) flag_l2_8;
  assign flag_l3_5 = flag_l2_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1726" *) flag_l2_10;
  assign flag_l3_6 = flag_l2_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1727" *) flag_l2_12;
  assign flag_l3_7 = flag_l2_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1728" *) flag_l2_14;
  assign flag_l3_8 = flag_l2_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1729" *) flag_l2_16;
  assign flag_l3_9 = flag_l2_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1730" *) flag_l2_18;
  assign flag_l3_10 = flag_l2_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1731" *) flag_l2_20;
  assign flag_l3_11 = flag_l2_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1732" *) flag_l2_22;
  assign flag_l3_12 = flag_l2_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1733" *) flag_l2_24;
  assign flag_l3_13 = flag_l2_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1734" *) flag_l2_26;
  assign flag_l3_14 = flag_l2_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1735" *) flag_l2_28;
  assign flag_l4_0 = flag_l3_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1736" *) flag_l3_0;
  assign flag_l4_1 = flag_l3_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1737" *) flag_l3_2;
  assign flag_l4_2 = flag_l3_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1738" *) flag_l3_4;
  assign flag_l4_3 = flag_l3_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1739" *) flag_l3_6;
  assign flag_l4_4 = flag_l3_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1740" *) flag_l3_8;
  assign flag_l4_5 = flag_l3_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1741" *) flag_l3_10;
  assign flag_l4_6 = flag_l3_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1742" *) flag_l3_12;
  assign flag_l5_0 = flag_l4_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1743" *) flag_l4_0;
  assign flag_l5_1 = flag_l4_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1744" *) flag_l4_2;
  assign flag_l5_2 = flag_l4_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1745" *) flag_l4_4;
  assign flag_l6_0 = flag_l5_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1746" *) flag_l5_0;
  assign _2479_ = cq_rd_credit[0] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2633" *) rd_take0;
  assign _2480_ = cq_rd_credit[1] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2729" *) rd_take1;
  assign _2481_ = cq_rd_credit[2] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2825" *) rd_take2;
  assign _2482_ = cq_rd_credit[3] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2921" *) rd_take3;
  assign _2483_ = cq_rd_credit[4] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3017" *) rd_take4;
  assign _2484_ = cq_rd_credit[5] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3113" *) rd_take5;
  assign _2485_ = cq_rd_credit[6] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3209" *) rd_take6;
  assign _2486_ = cq_rd_credit[7] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3305" *) rd_take7;
  assign _2487_ = cq_rd_credit[8] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3401" *) rd_take8;
  assign _2488_ = cq_rd_credit[9] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3497" *) rd_take9;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_take_thread_id_last <= 4'b0000;
    else
      cq_rd_take_thread_id_last <= _0031_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd9_credits <= 9'b000000000;
    else
      cq_rd9_credits <= _0018_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd9_credits_ne0 <= 1'b0;
    else
      cq_rd9_credits_ne0 <= _0019_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid9_0_vld <= 1'b0;
    else
      rd_skid9_0_vld <= _0101_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid9_1_vld <= 1'b0;
    else
      rd_skid9_1_vld <= _0103_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid9_2_vld <= 1'b0;
    else
      rd_skid9_2_vld <= _0105_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid9_0 <= _0100_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid9_1 <= _0102_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid9_2 <= _0104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd9_prdy_d <= 1'b1;
    else
      cq_rd9_prdy_d <= cq_rd9_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd8_credits <= 9'b000000000;
    else
      cq_rd8_credits <= _0016_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd8_credits_ne0 <= 1'b0;
    else
      cq_rd8_credits_ne0 <= _0017_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid8_0_vld <= 1'b0;
    else
      rd_skid8_0_vld <= _0095_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid8_1_vld <= 1'b0;
    else
      rd_skid8_1_vld <= _0097_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid8_2_vld <= 1'b0;
    else
      rd_skid8_2_vld <= _0099_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid8_0 <= _0094_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid8_1 <= _0096_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid8_2 <= _0098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd8_prdy_d <= 1'b1;
    else
      cq_rd8_prdy_d <= cq_rd8_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd7_credits <= 9'b000000000;
    else
      cq_rd7_credits <= _0014_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd7_credits_ne0 <= 1'b0;
    else
      cq_rd7_credits_ne0 <= _0015_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid7_0_vld <= 1'b0;
    else
      rd_skid7_0_vld <= _0089_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid7_1_vld <= 1'b0;
    else
      rd_skid7_1_vld <= _0091_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid7_2_vld <= 1'b0;
    else
      rd_skid7_2_vld <= _0093_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid7_0 <= _0088_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid7_1 <= _0090_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid7_2 <= _0092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd7_prdy_d <= 1'b1;
    else
      cq_rd7_prdy_d <= cq_rd7_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd6_credits <= 9'b000000000;
    else
      cq_rd6_credits <= _0012_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd6_credits_ne0 <= 1'b0;
    else
      cq_rd6_credits_ne0 <= _0013_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid6_0_vld <= 1'b0;
    else
      rd_skid6_0_vld <= _0083_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid6_1_vld <= 1'b0;
    else
      rd_skid6_1_vld <= _0085_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid6_2_vld <= 1'b0;
    else
      rd_skid6_2_vld <= _0087_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid6_0 <= _0082_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid6_1 <= _0084_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid6_2 <= _0086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd6_prdy_d <= 1'b1;
    else
      cq_rd6_prdy_d <= cq_rd6_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd5_credits <= 9'b000000000;
    else
      cq_rd5_credits <= _0010_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd5_credits_ne0 <= 1'b0;
    else
      cq_rd5_credits_ne0 <= _0011_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid5_0_vld <= 1'b0;
    else
      rd_skid5_0_vld <= _0077_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid5_1_vld <= 1'b0;
    else
      rd_skid5_1_vld <= _0079_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid5_2_vld <= 1'b0;
    else
      rd_skid5_2_vld <= _0081_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid5_0 <= _0076_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid5_1 <= _0078_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid5_2 <= _0080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd5_prdy_d <= 1'b1;
    else
      cq_rd5_prdy_d <= cq_rd5_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_credits <= 9'b000000000;
    else
      cq_rd4_credits <= _0008_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_credits_ne0 <= 1'b0;
    else
      cq_rd4_credits_ne0 <= _0009_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_0_vld <= 1'b0;
    else
      rd_skid4_0_vld <= _0071_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_1_vld <= 1'b0;
    else
      rd_skid4_1_vld <= _0073_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_2_vld <= 1'b0;
    else
      rd_skid4_2_vld <= _0075_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_0 <= _0070_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_1 <= _0072_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_2 <= _0074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_prdy_d <= 1'b1;
    else
      cq_rd4_prdy_d <= cq_rd4_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_credits <= 9'b000000000;
    else
      cq_rd3_credits <= _0006_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_credits_ne0 <= 1'b0;
    else
      cq_rd3_credits_ne0 <= _0007_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_0_vld <= 1'b0;
    else
      rd_skid3_0_vld <= _0065_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_1_vld <= 1'b0;
    else
      rd_skid3_1_vld <= _0067_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_2_vld <= 1'b0;
    else
      rd_skid3_2_vld <= _0069_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_0 <= _0064_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_1 <= _0066_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_2 <= _0068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_prdy_d <= 1'b1;
    else
      cq_rd3_prdy_d <= cq_rd3_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_credits <= 9'b000000000;
    else
      cq_rd2_credits <= _0004_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_credits_ne0 <= 1'b0;
    else
      cq_rd2_credits_ne0 <= _0005_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_0_vld <= 1'b0;
    else
      rd_skid2_0_vld <= _0059_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_1_vld <= 1'b0;
    else
      rd_skid2_1_vld <= _0061_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_2_vld <= 1'b0;
    else
      rd_skid2_2_vld <= _0063_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_0 <= _0058_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_1 <= _0060_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_2 <= _0062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_prdy_d <= 1'b1;
    else
      cq_rd2_prdy_d <= cq_rd2_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_credits <= 9'b000000000;
    else
      cq_rd1_credits <= _0002_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_credits_ne0 <= 1'b0;
    else
      cq_rd1_credits_ne0 <= _0003_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_0_vld <= 1'b0;
    else
      rd_skid1_0_vld <= _0053_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_1_vld <= 1'b0;
    else
      rd_skid1_1_vld <= _0055_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_2_vld <= 1'b0;
    else
      rd_skid1_2_vld <= _0057_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_0 <= _0052_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_1 <= _0054_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_2 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_prdy_d <= 1'b1;
    else
      cq_rd1_prdy_d <= cq_rd1_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_credits <= 9'b000000000;
    else
      cq_rd0_credits <= _0000_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_credits_ne0 <= 1'b0;
    else
      cq_rd0_credits_ne0 <= _0001_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_0_vld <= 1'b0;
    else
      rd_skid0_0_vld <= _0047_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_1_vld <= 1'b0;
    else
      rd_skid0_1_vld <= _0049_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_2_vld <= 1'b0;
    else
      rd_skid0_2_vld <= _0051_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_0 <= _0046_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_1 <= _0048_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_2 <= _0050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_prdy_d <= 1'b1;
    else
      cq_rd0_prdy_d <= cq_rd0_prdy;
  always @(posedge nvdla_core_clk_mgated)
      rd_adr_dly <= _0044_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_take_dly <= 1'b0;
    else
      rd_take_dly <= cq_rd_take;
  always @(posedge nvdla_core_clk_mgated)
      head0 <= _0034_;
  always @(posedge nvdla_core_clk_mgated)
      tail0 <= _0107_;
  always @(posedge nvdla_core_clk_mgated)
      head1 <= _0035_;
  always @(posedge nvdla_core_clk_mgated)
      tail1 <= _0108_;
  always @(posedge nvdla_core_clk_mgated)
      head2 <= _0036_;
  always @(posedge nvdla_core_clk_mgated)
      tail2 <= _0109_;
  always @(posedge nvdla_core_clk_mgated)
      head3 <= _0037_;
  always @(posedge nvdla_core_clk_mgated)
      tail3 <= _0110_;
  always @(posedge nvdla_core_clk_mgated)
      head4 <= _0038_;
  always @(posedge nvdla_core_clk_mgated)
      tail4 <= _0111_;
  always @(posedge nvdla_core_clk_mgated)
      head5 <= _0039_;
  always @(posedge nvdla_core_clk_mgated)
      tail5 <= _0112_;
  always @(posedge nvdla_core_clk_mgated)
      head6 <= _0040_;
  always @(posedge nvdla_core_clk_mgated)
      tail6 <= _0113_;
  always @(posedge nvdla_core_clk_mgated)
      head7 <= _0041_;
  always @(posedge nvdla_core_clk_mgated)
      tail7 <= _0114_;
  always @(posedge nvdla_core_clk_mgated)
      head8 <= _0042_;
  always @(posedge nvdla_core_clk_mgated)
      tail8 <= _0115_;
  always @(posedge nvdla_core_clk_mgated)
      head9 <= _0043_;
  always @(posedge nvdla_core_clk_mgated)
      tail9 <= _0116_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      update_head <= 10'b0000000000;
    else
      update_head <= _0117_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count0 <= 9'b000000000;
    else
      cq_rd_count0 <= _0020_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count1 <= 9'b000000000;
    else
      cq_rd_count1 <= _0021_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count2 <= 9'b000000000;
    else
      cq_rd_count2 <= _0022_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count3 <= 9'b000000000;
    else
      cq_rd_count3 <= _0023_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count4 <= 9'b000000000;
    else
      cq_rd_count4 <= _0024_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count5 <= 9'b000000000;
    else
      cq_rd_count5 <= _0025_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count6 <= 9'b000000000;
    else
      cq_rd_count6 <= _0026_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count7 <= 9'b000000000;
    else
      cq_rd_count7 <= _0027_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count8 <= 9'b000000000;
    else
      cq_rd_count8 <= _0028_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count9 <= 9'b000000000;
    else
      cq_rd_count9 <= _0029_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_take_n_dly <= 10'b0000000000;
    else
      rd_take_n_dly <= _0106_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_credit <= 10'b0000000000;
    else
      cq_rd_credit <= _0030_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pushing_q <= 1'b0;
    else
      rd_pushing_q <= _0045_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      free_adr_mask <= 255'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    else
      free_adr_mask <= _0033_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_wr_busy_int <= 1'b0;
    else
      cq_wr_busy_int <= cq_wr_busy_next;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_wr_count <= 9'b000000000;
    else
      cq_wr_count <= _0032_;
  assign _0031_ = cq_rd_take ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3619" *) cq_rd_take_thread_id : cq_rd_take_thread_id_last;
  assign _0019_ = _2488_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3497" *) _2600_ : cq_rd9_credits_ne0;
  assign _0018_ = _2488_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3497" *) cq_rd9_credits_next : cq_rd9_credits;
  assign _0104_ = _1461_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3457" *) _2599_ : rd_skid9_2;
  assign _2489_ = _1458_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3447" *) rd_skid9_2 : rd_skid9_1;
  assign _0102_ = _1457_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3445" *) _2599_ : _2489_;
  assign _2490_ = _1454_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3435" *) rd_skid9_1 : rd_skid9_0;
  assign _0100_ = _1453_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3433" *) _2598_ : _2490_;
  assign _0017_ = _2487_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3401" *) _2597_ : cq_rd8_credits_ne0;
  assign _0016_ = _2487_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3401" *) cq_rd8_credits_next : cq_rd8_credits;
  assign _0098_ = _1438_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3361" *) _2596_ : rd_skid8_2;
  assign _2491_ = _1434_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3351" *) rd_skid8_2 : rd_skid8_1;
  assign _0096_ = _1433_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3349" *) _2596_ : _2491_;
  assign _2492_ = _1430_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3339" *) rd_skid8_1 : rd_skid8_0;
  assign _0094_ = _1429_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3337" *) _2595_ : _2492_;
  assign _0015_ = _2486_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3305" *) _2594_ : cq_rd7_credits_ne0;
  assign _0014_ = _2486_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3305" *) cq_rd7_credits_next : cq_rd7_credits;
  assign _0092_ = _1414_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3265" *) _2593_ : rd_skid7_2;
  assign _2493_ = _1410_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3255" *) rd_skid7_2 : rd_skid7_1;
  assign _0090_ = _1409_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3253" *) _2593_ : _2493_;
  assign _2494_ = _1407_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3243" *) rd_skid7_1 : rd_skid7_0;
  assign _0088_ = _1406_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3241" *) _2592_ : _2494_;
  assign _0013_ = _2485_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3209" *) _2591_ : cq_rd6_credits_ne0;
  assign _0012_ = _2485_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3209" *) cq_rd6_credits_next : cq_rd6_credits;
  assign _0086_ = _1390_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3169" *) _2590_ : rd_skid6_2;
  assign _2495_ = _1386_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3159" *) rd_skid6_2 : rd_skid6_1;
  assign _0084_ = _1385_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3157" *) _2590_ : _2495_;
  assign _2496_ = _1383_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3147" *) rd_skid6_1 : rd_skid6_0;
  assign _0082_ = _1382_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3145" *) _2589_ : _2496_;
  assign _0011_ = _2484_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3113" *) _2588_ : cq_rd5_credits_ne0;
  assign _0010_ = _2484_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3113" *) cq_rd5_credits_next : cq_rd5_credits;
  assign _0080_ = _1366_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3073" *) _2587_ : rd_skid5_2;
  assign _2497_ = _1363_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3063" *) rd_skid5_2 : rd_skid5_1;
  assign _0078_ = _1362_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3061" *) _2587_ : _2497_;
  assign _2498_ = _1359_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3051" *) rd_skid5_1 : rd_skid5_0;
  assign _0076_ = _1358_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3049" *) _2586_ : _2498_;
  assign _0009_ = _2483_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3017" *) _2585_ : cq_rd4_credits_ne0;
  assign _0008_ = _2483_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3017" *) cq_rd4_credits_next : cq_rd4_credits;
  assign _0074_ = _1342_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2977" *) _2584_ : rd_skid4_2;
  assign _2499_ = _1339_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2967" *) rd_skid4_2 : rd_skid4_1;
  assign _0072_ = _1338_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2965" *) _2584_ : _2499_;
  assign _2500_ = _1335_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2955" *) rd_skid4_1 : rd_skid4_0;
  assign _0070_ = _1334_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2953" *) _2583_ : _2500_;
  assign _0007_ = _2482_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2921" *) _2582_ : cq_rd3_credits_ne0;
  assign _0006_ = _2482_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2921" *) cq_rd3_credits_next : cq_rd3_credits;
  assign _0068_ = _1318_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2881" *) _2581_ : rd_skid3_2;
  assign _2501_ = _1315_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2871" *) rd_skid3_2 : rd_skid3_1;
  assign _0066_ = _1314_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2869" *) _2581_ : _2501_;
  assign _2502_ = _1311_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2859" *) rd_skid3_1 : rd_skid3_0;
  assign _0064_ = _1310_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2857" *) _2580_ : _2502_;
  assign _0005_ = _2481_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2825" *) _2579_ : cq_rd2_credits_ne0;
  assign _0004_ = _2481_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2825" *) cq_rd2_credits_next : cq_rd2_credits;
  assign _0062_ = _1294_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2785" *) _2578_ : rd_skid2_2;
  assign _2503_ = _1291_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2775" *) rd_skid2_2 : rd_skid2_1;
  assign _0060_ = _1290_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2773" *) _2578_ : _2503_;
  assign _2504_ = _1288_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2763" *) rd_skid2_1 : rd_skid2_0;
  assign _0058_ = _1287_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2761" *) _2577_ : _2504_;
  assign _0003_ = _2480_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2729" *) _2576_ : cq_rd1_credits_ne0;
  assign _0002_ = _2480_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2729" *) cq_rd1_credits_next : cq_rd1_credits;
  assign _0056_ = _1270_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2689" *) _2575_ : rd_skid1_2;
  assign _2505_ = _1267_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2679" *) rd_skid1_2 : rd_skid1_1;
  assign _0054_ = _1266_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2677" *) _2575_ : _2505_;
  assign _2506_ = _1264_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2667" *) rd_skid1_1 : rd_skid1_0;
  assign _0052_ = _1263_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2665" *) _2574_ : _2506_;
  assign _0001_ = _2479_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2633" *) _2573_ : cq_rd0_credits_ne0;
  assign _0000_ = _2479_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2633" *) cq_rd0_credits_next : cq_rd0_credits;
  assign _0050_ = _1247_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2593" *) _2572_ : rd_skid0_2;
  assign _2507_ = _1243_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2583" *) rd_skid0_2 : rd_skid0_1;
  assign _0048_ = _1242_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2581" *) _2572_ : _2507_;
  assign _2508_ = _1240_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2571" *) rd_skid0_1 : rd_skid0_0;
  assign _0046_ = _1239_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2569" *) _2571_ : _2508_;
  assign _0044_ = cq_rd_take ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2538" *) adr_ram_rd_adr : rd_adr_dly;
  function [7:0] _5599_;
    input [7:0] a;
    input [79:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2517|./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2507" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _5599_ = b[7:0];
      10'b????????1?:
        _5599_ = b[15:8];
      10'b???????1??:
        _5599_ = b[23:16];
      10'b??????1???:
        _5599_ = b[31:24];
      10'b?????1????:
        _5599_ = b[39:32];
      10'b????1?????:
        _5599_ = b[47:40];
      10'b???1??????:
        _5599_ = b[55:48];
      10'b??1???????:
        _5599_ = b[63:56];
      10'b?1????????:
        _5599_ = b[71:64];
      10'b1?????????:
        _5599_ = b[79:72];
      default:
        _5599_ = a;
    endcase
  endfunction
  assign adr_ram_rd_adr = _5599_(8'b00000000, { _2561_, _2562_, _2563_, _2564_, _2565_, _2566_, _2567_, _2568_, _2569_, _2570_ }, { _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_ });
  function [0:0] _5600_;
    input [0:0] a;
    input [9:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2483|./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2473" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _5600_ = b[0:0];
      10'b????????1?:
        _5600_ = b[1:1];
      10'b???????1??:
        _5600_ = b[2:2];
      10'b??????1???:
        _5600_ = b[3:3];
      10'b?????1????:
        _5600_ = b[4:4];
      10'b????1?????:
        _5600_ = b[5:5];
      10'b???1??????:
        _5600_ = b[6:6];
      10'b??1???????:
        _5600_ = b[7:7];
      10'b?1????????:
        _5600_ = b[8:8];
      10'b1?????????:
        _5600_ = b[9:9];
      default:
        _5600_ = a;
    endcase
  endfunction
  assign adr_ram_rd_enable = _5600_(1'b0, { _1213_, _1214_, _1215_, _1216_, _1217_, _1218_, _1219_, _1220_, _1221_, _1222_ }, { _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_ });
  function [0:0] _5601_;
    input [0:0] a;
    input [9:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2466|./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2456" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _5601_ = b[0:0];
      10'b????????1?:
        _5601_ = b[1:1];
      10'b???????1??:
        _5601_ = b[2:2];
      10'b??????1???:
        _5601_ = b[3:3];
      10'b?????1????:
        _5601_ = b[4:4];
      10'b????1?????:
        _5601_ = b[5:5];
      10'b???1??????:
        _5601_ = b[6:6];
      10'b??1???????:
        _5601_ = b[7:7];
      10'b?1????????:
        _5601_ = b[8:8];
      10'b1?????????:
        _5601_ = b[9:9];
      default:
        _5601_ = a;
    endcase
  endfunction
  assign adr_ram_wr_enable = _5601_(1'b0, { _1202_, _1203_, _1204_, _1206_, _1207_, _1208_, _1209_, _1210_, _1211_, _1212_ }, { _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_ });
  function [7:0] _5602_;
    input [7:0] a;
    input [79:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2449|./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2439" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _5602_ = b[7:0];
      10'b????????1?:
        _5602_ = b[15:8];
      10'b???????1??:
        _5602_ = b[23:16];
      10'b??????1???:
        _5602_ = b[31:24];
      10'b?????1????:
        _5602_ = b[39:32];
      10'b????1?????:
        _5602_ = b[47:40];
      10'b???1??????:
        _5602_ = b[55:48];
      10'b??1???????:
        _5602_ = b[63:56];
      10'b?1????????:
        _5602_ = b[71:64];
      10'b1?????????:
        _5602_ = b[79:72];
      default:
        _5602_ = a;
    endcase
  endfunction
  assign adr_ram_wr_adr = _5602_(8'b00000000, { tail0, tail1, tail2, tail3, tail4, tail5, tail6, tail7, tail8, tail9 }, { _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_ });
  assign _0116_ = rd_pushing9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2411" *) adr_ram_wr_data : tail9;
  assign _2509_ = update_head[9] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2423" *) adr_ram_rd_data : head9;
  assign _0043_ = _2242_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2421" *) adr_ram_wr_data : _2509_;
  assign _0115_ = rd_pushing8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2396" *) adr_ram_wr_data : tail8;
  assign _2510_ = update_head[8] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2408" *) adr_ram_rd_data : head8;
  assign _0042_ = _2241_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2406" *) adr_ram_wr_data : _2510_;
  assign _0114_ = rd_pushing7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2381" *) adr_ram_wr_data : tail7;
  assign _2511_ = update_head[7] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2393" *) adr_ram_rd_data : head7;
  assign _0041_ = _2240_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2391" *) adr_ram_wr_data : _2511_;
  assign _0113_ = rd_pushing6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2366" *) adr_ram_wr_data : tail6;
  assign _2512_ = update_head[6] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2378" *) adr_ram_rd_data : head6;
  assign _0040_ = _2239_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2376" *) adr_ram_wr_data : _2512_;
  assign _0112_ = rd_pushing5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2351" *) adr_ram_wr_data : tail5;
  assign _2513_ = update_head[5] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2363" *) adr_ram_rd_data : head5;
  assign _0039_ = _2238_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2361" *) adr_ram_wr_data : _2513_;
  assign _0111_ = rd_pushing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2336" *) adr_ram_wr_data : tail4;
  assign _2514_ = update_head[4] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2348" *) adr_ram_rd_data : head4;
  assign _0038_ = _2237_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2346" *) adr_ram_wr_data : _2514_;
  assign _0110_ = rd_pushing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2321" *) adr_ram_wr_data : tail3;
  assign _2515_ = update_head[3] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2333" *) adr_ram_rd_data : head3;
  assign _0037_ = _2236_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2331" *) adr_ram_wr_data : _2515_;
  assign _0109_ = rd_pushing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2306" *) adr_ram_wr_data : tail2;
  assign _2516_ = update_head[2] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2318" *) adr_ram_rd_data : head2;
  assign _0036_ = _2235_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2316" *) adr_ram_wr_data : _2516_;
  assign _0108_ = rd_pushing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2291" *) adr_ram_wr_data : tail1;
  assign _2517_ = update_head[1] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2303" *) adr_ram_rd_data : head1;
  assign _0035_ = _2234_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2301" *) adr_ram_wr_data : _2517_;
  assign _0107_ = rd_pushing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2276" *) adr_ram_wr_data : tail0;
  assign _2518_ = update_head[0] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2288" *) adr_ram_rd_data : head0;
  assign _0034_ = _2233_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2286" *) adr_ram_wr_data : _2518_;
  assign _0117_ = _2232_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2264" *) update_head_next : update_head;
  assign _0029_ = _2519_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2237" *) rd_count9_next : cq_rd_count9;
  assign _0028_ = _2520_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2228" *) rd_count8_next : cq_rd_count8;
  assign _0027_ = _2521_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2219" *) rd_count7_next : cq_rd_count7;
  assign _0026_ = _2522_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2210" *) rd_count6_next : cq_rd_count6;
  assign _0025_ = _2523_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2201" *) rd_count5_next : cq_rd_count5;
  assign _0024_ = _2524_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2192" *) rd_count4_next : cq_rd_count4;
  assign _0023_ = _2525_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2183" *) rd_count3_next : cq_rd_count3;
  assign _0022_ = _2526_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2174" *) rd_count2_next : cq_rd_count2;
  assign _0021_ = _2527_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2165" *) rd_count1_next : cq_rd_count1;
  assign _0020_ = _2528_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2156" *) rd_count0_next : cq_rd_count0;
  assign _0106_ = update_rd_take_n_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2076" *) { rd_take9, rd_take8, rd_take7, rd_take6, rd_take5, rd_take4, rd_take3, rd_take2, rd_take1, rd_take0 } : rd_take_n_dly;
  assign _0030_[9] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing9 : cq_rd_credit[9];
  assign _0030_[8] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing8 : cq_rd_credit[8];
  assign _0030_[7] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing7 : cq_rd_credit[7];
  assign _0030_[6] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing6 : cq_rd_credit[6];
  assign _0030_[5] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing5 : cq_rd_credit[5];
  assign _0030_[4] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing4 : cq_rd_credit[4];
  assign _0030_[3] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing3 : cq_rd_credit[3];
  assign _0030_[2] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing2 : cq_rd_credit[2];
  assign _0030_[1] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing1 : cq_rd_credit[1];
  assign _0030_[0] = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing0 : cq_rd_credit[0];
  assign _0045_ = _2230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2012" *) rd_pushing : rd_pushing_q;
  assign _0346_ = _1162_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1496" *) 1'b0 : free_adr_mask[254];
  assign free_adr_mask_next[254] = _1161_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1494" *) 1'b1 : _0346_;
  assign _0344_ = _1160_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1491" *) 1'b0 : free_adr_mask[253];
  assign free_adr_mask_next[253] = _1159_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1489" *) 1'b1 : _0344_;
  assign _0343_ = _1158_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1486" *) 1'b0 : free_adr_mask[252];
  assign free_adr_mask_next[252] = _1157_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1484" *) 1'b1 : _0343_;
  assign _0342_ = _1156_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1481" *) 1'b0 : free_adr_mask[251];
  assign free_adr_mask_next[251] = _1155_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1479" *) 1'b1 : _0342_;
  assign _0341_ = _1154_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1476" *) 1'b0 : free_adr_mask[250];
  assign free_adr_mask_next[250] = _1153_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1474" *) 1'b1 : _0341_;
  assign _0340_ = _1152_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1471" *) 1'b0 : free_adr_mask[249];
  assign free_adr_mask_next[249] = _1151_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1469" *) 1'b1 : _0340_;
  assign _0338_ = _1150_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1466" *) 1'b0 : free_adr_mask[248];
  assign free_adr_mask_next[248] = _1149_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1464" *) 1'b1 : _0338_;
  assign _0337_ = _1148_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1461" *) 1'b0 : free_adr_mask[247];
  assign free_adr_mask_next[247] = _1147_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1459" *) 1'b1 : _0337_;
  assign _0336_ = _1146_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1456" *) 1'b0 : free_adr_mask[246];
  assign free_adr_mask_next[246] = _1145_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1454" *) 1'b1 : _0336_;
  assign _0335_ = _1144_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1451" *) 1'b0 : free_adr_mask[245];
  assign free_adr_mask_next[245] = _1143_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1449" *) 1'b1 : _0335_;
  assign _0334_ = _1142_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1446" *) 1'b0 : free_adr_mask[244];
  assign free_adr_mask_next[244] = _1141_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1444" *) 1'b1 : _0334_;
  assign _0332_ = _1140_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1441" *) 1'b0 : free_adr_mask[243];
  assign free_adr_mask_next[243] = _1139_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1439" *) 1'b1 : _0332_;
  assign _0331_ = _1138_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1436" *) 1'b0 : free_adr_mask[242];
  assign free_adr_mask_next[242] = _1137_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1434" *) 1'b1 : _0331_;
  assign _0330_ = _1136_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1431" *) 1'b0 : free_adr_mask[241];
  assign free_adr_mask_next[241] = _1135_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1429" *) 1'b1 : _0330_;
  assign _0329_ = _1134_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1426" *) 1'b0 : free_adr_mask[240];
  assign free_adr_mask_next[240] = _1133_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1424" *) 1'b1 : _0329_;
  assign _0328_ = _1132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1421" *) 1'b0 : free_adr_mask[239];
  assign free_adr_mask_next[239] = _1131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1419" *) 1'b1 : _0328_;
  assign _0327_ = _1130_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1416" *) 1'b0 : free_adr_mask[238];
  assign free_adr_mask_next[238] = _1129_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1414" *) 1'b1 : _0327_;
  assign _0326_ = _1128_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1411" *) 1'b0 : free_adr_mask[237];
  assign free_adr_mask_next[237] = _1127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1409" *) 1'b1 : _0326_;
  assign _0325_ = _1126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1406" *) 1'b0 : free_adr_mask[236];
  assign free_adr_mask_next[236] = _1125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1404" *) 1'b1 : _0325_;
  assign _0324_ = _1124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1401" *) 1'b0 : free_adr_mask[235];
  assign free_adr_mask_next[235] = _1123_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1399" *) 1'b1 : _0324_;
  assign _0323_ = _1122_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1396" *) 1'b0 : free_adr_mask[234];
  assign free_adr_mask_next[234] = _1121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1394" *) 1'b1 : _0323_;
  assign _0321_ = _1120_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1391" *) 1'b0 : free_adr_mask[233];
  assign free_adr_mask_next[233] = _1119_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1389" *) 1'b1 : _0321_;
  assign _0320_ = _1118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1386" *) 1'b0 : free_adr_mask[232];
  assign free_adr_mask_next[232] = _1117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1384" *) 1'b1 : _0320_;
  assign _0319_ = _1116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1381" *) 1'b0 : free_adr_mask[231];
  assign free_adr_mask_next[231] = _1115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1379" *) 1'b1 : _0319_;
  assign _0318_ = _1114_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1376" *) 1'b0 : free_adr_mask[230];
  assign free_adr_mask_next[230] = _1113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1374" *) 1'b1 : _0318_;
  assign _0317_ = _1112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1371" *) 1'b0 : free_adr_mask[229];
  assign free_adr_mask_next[229] = _1111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1369" *) 1'b1 : _0317_;
  assign _0316_ = _1110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1366" *) 1'b0 : free_adr_mask[228];
  assign free_adr_mask_next[228] = _1109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1364" *) 1'b1 : _0316_;
  assign _0315_ = _1108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1361" *) 1'b0 : free_adr_mask[227];
  assign free_adr_mask_next[227] = _1107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1359" *) 1'b1 : _0315_;
  assign _0314_ = _1106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1356" *) 1'b0 : free_adr_mask[226];
  assign free_adr_mask_next[226] = _1105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1354" *) 1'b1 : _0314_;
  assign _0313_ = _1104_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1351" *) 1'b0 : free_adr_mask[225];
  assign free_adr_mask_next[225] = _1103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1349" *) 1'b1 : _0313_;
  assign _0312_ = _1102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1346" *) 1'b0 : free_adr_mask[224];
  assign free_adr_mask_next[224] = _1101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1344" *) 1'b1 : _0312_;
  assign _0310_ = _1100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1341" *) 1'b0 : free_adr_mask[223];
  assign free_adr_mask_next[223] = _1099_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1339" *) 1'b1 : _0310_;
  assign _0309_ = _1098_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1336" *) 1'b0 : free_adr_mask[222];
  assign free_adr_mask_next[222] = _1097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1334" *) 1'b1 : _0309_;
  assign _0308_ = _1096_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1331" *) 1'b0 : free_adr_mask[221];
  assign free_adr_mask_next[221] = _1095_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1329" *) 1'b1 : _0308_;
  assign _0307_ = _1094_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1326" *) 1'b0 : free_adr_mask[220];
  assign free_adr_mask_next[220] = _1093_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1324" *) 1'b1 : _0307_;
  assign _0306_ = _1092_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1321" *) 1'b0 : free_adr_mask[219];
  assign free_adr_mask_next[219] = _1091_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1319" *) 1'b1 : _0306_;
  assign _0305_ = _1090_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1316" *) 1'b0 : free_adr_mask[218];
  assign free_adr_mask_next[218] = _1089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1314" *) 1'b1 : _0305_;
  assign _0304_ = _1088_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1311" *) 1'b0 : free_adr_mask[217];
  assign free_adr_mask_next[217] = _1087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1309" *) 1'b1 : _0304_;
  assign _0303_ = _1086_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1306" *) 1'b0 : free_adr_mask[216];
  assign free_adr_mask_next[216] = _1085_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1304" *) 1'b1 : _0303_;
  assign _0302_ = _1084_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1301" *) 1'b0 : free_adr_mask[215];
  assign free_adr_mask_next[215] = _1083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1299" *) 1'b1 : _0302_;
  assign _0301_ = _1082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1296" *) 1'b0 : free_adr_mask[214];
  assign free_adr_mask_next[214] = _1081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1294" *) 1'b1 : _0301_;
  assign _0299_ = _1080_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1291" *) 1'b0 : free_adr_mask[213];
  assign free_adr_mask_next[213] = _1079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1289" *) 1'b1 : _0299_;
  assign _0298_ = _1078_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1286" *) 1'b0 : free_adr_mask[212];
  assign free_adr_mask_next[212] = _1077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1284" *) 1'b1 : _0298_;
  assign _0297_ = _1076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1281" *) 1'b0 : free_adr_mask[211];
  assign free_adr_mask_next[211] = _1075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1279" *) 1'b1 : _0297_;
  assign _0296_ = _1074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1276" *) 1'b0 : free_adr_mask[210];
  assign free_adr_mask_next[210] = _1073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1274" *) 1'b1 : _0296_;
  assign _0295_ = _1072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1271" *) 1'b0 : free_adr_mask[209];
  assign free_adr_mask_next[209] = _1071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1269" *) 1'b1 : _0295_;
  assign _0294_ = _1070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1266" *) 1'b0 : free_adr_mask[208];
  assign free_adr_mask_next[208] = _1069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1264" *) 1'b1 : _0294_;
  assign _0293_ = _1068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1261" *) 1'b0 : free_adr_mask[207];
  assign free_adr_mask_next[207] = _1067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1259" *) 1'b1 : _0293_;
  assign _0292_ = _1066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1256" *) 1'b0 : free_adr_mask[206];
  assign free_adr_mask_next[206] = _1065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1254" *) 1'b1 : _0292_;
  assign _0291_ = _1064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1251" *) 1'b0 : free_adr_mask[205];
  assign free_adr_mask_next[205] = _1063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1249" *) 1'b1 : _0291_;
  assign _0290_ = _1062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1246" *) 1'b0 : free_adr_mask[204];
  assign free_adr_mask_next[204] = _1061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1244" *) 1'b1 : _0290_;
  assign _0288_ = _1060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1241" *) 1'b0 : free_adr_mask[203];
  assign free_adr_mask_next[203] = _1059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1239" *) 1'b1 : _0288_;
  assign _0287_ = _1058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1236" *) 1'b0 : free_adr_mask[202];
  assign free_adr_mask_next[202] = _1057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1234" *) 1'b1 : _0287_;
  assign _0286_ = _1056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1231" *) 1'b0 : free_adr_mask[201];
  assign free_adr_mask_next[201] = _1055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1229" *) 1'b1 : _0286_;
  assign _0285_ = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1226" *) 1'b0 : free_adr_mask[200];
  assign free_adr_mask_next[200] = _1053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1224" *) 1'b1 : _0285_;
  assign _0284_ = _1052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1221" *) 1'b0 : free_adr_mask[199];
  assign free_adr_mask_next[199] = _1051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1219" *) 1'b1 : _0284_;
  assign _0283_ = _1050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1216" *) 1'b0 : free_adr_mask[198];
  assign free_adr_mask_next[198] = _1049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1214" *) 1'b1 : _0283_;
  assign _0282_ = _1048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1211" *) 1'b0 : free_adr_mask[197];
  assign free_adr_mask_next[197] = _1047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1209" *) 1'b1 : _0282_;
  assign _0281_ = _1046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1206" *) 1'b0 : free_adr_mask[196];
  assign free_adr_mask_next[196] = _1045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1204" *) 1'b1 : _0281_;
  assign _0280_ = _1044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1201" *) 1'b0 : free_adr_mask[195];
  assign free_adr_mask_next[195] = _1043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1199" *) 1'b1 : _0280_;
  assign _0279_ = _1042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1196" *) 1'b0 : free_adr_mask[194];
  assign free_adr_mask_next[194] = _1041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1194" *) 1'b1 : _0279_;
  assign _0277_ = _1040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1191" *) 1'b0 : free_adr_mask[193];
  assign free_adr_mask_next[193] = _1039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1189" *) 1'b1 : _0277_;
  assign _0276_ = _1038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1186" *) 1'b0 : free_adr_mask[192];
  assign free_adr_mask_next[192] = _1037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1184" *) 1'b1 : _0276_;
  assign _0275_ = _1036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1181" *) 1'b0 : free_adr_mask[191];
  assign free_adr_mask_next[191] = _1035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1179" *) 1'b1 : _0275_;
  assign _0274_ = _1034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1176" *) 1'b0 : free_adr_mask[190];
  assign free_adr_mask_next[190] = _1033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1174" *) 1'b1 : _0274_;
  assign _0273_ = _1032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1171" *) 1'b0 : free_adr_mask[189];
  assign free_adr_mask_next[189] = _1031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1169" *) 1'b1 : _0273_;
  assign _0272_ = _1030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1166" *) 1'b0 : free_adr_mask[188];
  assign free_adr_mask_next[188] = _1029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1164" *) 1'b1 : _0272_;
  assign _0271_ = _1028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1161" *) 1'b0 : free_adr_mask[187];
  assign free_adr_mask_next[187] = _1027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1159" *) 1'b1 : _0271_;
  assign _0270_ = _1026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1156" *) 1'b0 : free_adr_mask[186];
  assign free_adr_mask_next[186] = _1025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1154" *) 1'b1 : _0270_;
  assign _0269_ = _1024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1151" *) 1'b0 : free_adr_mask[185];
  assign free_adr_mask_next[185] = _1023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1149" *) 1'b1 : _0269_;
  assign _0268_ = _1022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1146" *) 1'b0 : free_adr_mask[184];
  assign free_adr_mask_next[184] = _1021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1144" *) 1'b1 : _0268_;
  assign _0266_ = _1020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1141" *) 1'b0 : free_adr_mask[183];
  assign free_adr_mask_next[183] = _1019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1139" *) 1'b1 : _0266_;
  assign _0265_ = _1018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1136" *) 1'b0 : free_adr_mask[182];
  assign free_adr_mask_next[182] = _1017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1134" *) 1'b1 : _0265_;
  assign _0264_ = _1016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1131" *) 1'b0 : free_adr_mask[181];
  assign free_adr_mask_next[181] = _1015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1129" *) 1'b1 : _0264_;
  assign _0263_ = _1014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1126" *) 1'b0 : free_adr_mask[180];
  assign free_adr_mask_next[180] = _1013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1124" *) 1'b1 : _0263_;
  assign _0262_ = _1012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1121" *) 1'b0 : free_adr_mask[179];
  assign free_adr_mask_next[179] = _1011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1119" *) 1'b1 : _0262_;
  assign _0261_ = _1010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1116" *) 1'b0 : free_adr_mask[178];
  assign free_adr_mask_next[178] = _1009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1114" *) 1'b1 : _0261_;
  assign _0260_ = _1008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1111" *) 1'b0 : free_adr_mask[177];
  assign free_adr_mask_next[177] = _1007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1109" *) 1'b1 : _0260_;
  assign _0259_ = _1006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1106" *) 1'b0 : free_adr_mask[176];
  assign free_adr_mask_next[176] = _1005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1104" *) 1'b1 : _0259_;
  assign _0258_ = _1004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1101" *) 1'b0 : free_adr_mask[175];
  assign free_adr_mask_next[175] = _1003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1099" *) 1'b1 : _0258_;
  assign _0257_ = _1002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1096" *) 1'b0 : free_adr_mask[174];
  assign free_adr_mask_next[174] = _1001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1094" *) 1'b1 : _0257_;
  assign _0255_ = _1000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1091" *) 1'b0 : free_adr_mask[173];
  assign free_adr_mask_next[173] = _0999_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1089" *) 1'b1 : _0255_;
  assign _0254_ = _0998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1086" *) 1'b0 : free_adr_mask[172];
  assign free_adr_mask_next[172] = _0997_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1084" *) 1'b1 : _0254_;
  assign _0253_ = _0996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1081" *) 1'b0 : free_adr_mask[171];
  assign free_adr_mask_next[171] = _0995_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1079" *) 1'b1 : _0253_;
  assign _0252_ = _0994_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1076" *) 1'b0 : free_adr_mask[170];
  assign free_adr_mask_next[170] = _0993_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1074" *) 1'b1 : _0252_;
  assign _0251_ = _0992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1071" *) 1'b0 : free_adr_mask[169];
  assign free_adr_mask_next[169] = _0991_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1069" *) 1'b1 : _0251_;
  assign _0250_ = _0990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1066" *) 1'b0 : free_adr_mask[168];
  assign free_adr_mask_next[168] = _0989_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1064" *) 1'b1 : _0250_;
  assign _0249_ = _0988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1061" *) 1'b0 : free_adr_mask[167];
  assign free_adr_mask_next[167] = _0987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1059" *) 1'b1 : _0249_;
  assign _0248_ = _0986_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1056" *) 1'b0 : free_adr_mask[166];
  assign free_adr_mask_next[166] = _0985_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1054" *) 1'b1 : _0248_;
  assign _0247_ = _0984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1051" *) 1'b0 : free_adr_mask[165];
  assign free_adr_mask_next[165] = _0983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1049" *) 1'b1 : _0247_;
  assign _0246_ = _0982_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1046" *) 1'b0 : free_adr_mask[164];
  assign free_adr_mask_next[164] = _0981_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1044" *) 1'b1 : _0246_;
  assign _0244_ = _0980_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1041" *) 1'b0 : free_adr_mask[163];
  assign free_adr_mask_next[163] = _0979_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1039" *) 1'b1 : _0244_;
  assign _0243_ = _0978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1036" *) 1'b0 : free_adr_mask[162];
  assign free_adr_mask_next[162] = _0977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1034" *) 1'b1 : _0243_;
  assign _0242_ = _0976_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1031" *) 1'b0 : free_adr_mask[161];
  assign free_adr_mask_next[161] = _0975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1029" *) 1'b1 : _0242_;
  assign _0241_ = _0974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1026" *) 1'b0 : free_adr_mask[160];
  assign free_adr_mask_next[160] = _0973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1024" *) 1'b1 : _0241_;
  assign _0240_ = _0972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1021" *) 1'b0 : free_adr_mask[159];
  assign free_adr_mask_next[159] = _0971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1019" *) 1'b1 : _0240_;
  assign _0239_ = _0970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1016" *) 1'b0 : free_adr_mask[158];
  assign free_adr_mask_next[158] = _0969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1014" *) 1'b1 : _0239_;
  assign _0238_ = _0968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1011" *) 1'b0 : free_adr_mask[157];
  assign free_adr_mask_next[157] = _0967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1009" *) 1'b1 : _0238_;
  assign _0237_ = _0966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1006" *) 1'b0 : free_adr_mask[156];
  assign free_adr_mask_next[156] = _0965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1004" *) 1'b1 : _0237_;
  assign _0236_ = _0964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1001" *) 1'b0 : free_adr_mask[155];
  assign free_adr_mask_next[155] = _2138_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:999" *) 1'b1 : _0236_;
  assign _0235_ = _2137_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:996" *) 1'b0 : free_adr_mask[154];
  assign free_adr_mask_next[154] = _2136_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:994" *) 1'b1 : _0235_;
  assign _0233_ = _2135_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:991" *) 1'b0 : free_adr_mask[153];
  assign free_adr_mask_next[153] = _2134_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:989" *) 1'b1 : _0233_;
  assign _0232_ = _2133_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:986" *) 1'b0 : free_adr_mask[152];
  assign free_adr_mask_next[152] = _2132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:984" *) 1'b1 : _0232_;
  assign _0231_ = _2131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:981" *) 1'b0 : free_adr_mask[151];
  assign free_adr_mask_next[151] = _2130_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:979" *) 1'b1 : _0231_;
  assign _0230_ = _2129_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:976" *) 1'b0 : free_adr_mask[150];
  assign free_adr_mask_next[150] = _2128_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:974" *) 1'b1 : _0230_;
  assign _0229_ = _2127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:971" *) 1'b0 : free_adr_mask[149];
  assign free_adr_mask_next[149] = _2126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:969" *) 1'b1 : _0229_;
  assign _0227_ = _2125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:966" *) 1'b0 : free_adr_mask[148];
  assign free_adr_mask_next[148] = _2124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:964" *) 1'b1 : _0227_;
  assign _0226_ = _2123_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:961" *) 1'b0 : free_adr_mask[147];
  assign free_adr_mask_next[147] = _2122_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:959" *) 1'b1 : _0226_;
  assign _0225_ = _2121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:956" *) 1'b0 : free_adr_mask[146];
  assign free_adr_mask_next[146] = _2120_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:954" *) 1'b1 : _0225_;
  assign _0224_ = _2119_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:951" *) 1'b0 : free_adr_mask[145];
  assign free_adr_mask_next[145] = _2118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:949" *) 1'b1 : _0224_;
  assign _0223_ = _2117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:946" *) 1'b0 : free_adr_mask[144];
  assign free_adr_mask_next[144] = _2116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:944" *) 1'b1 : _0223_;
  assign _0221_ = _2115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:941" *) 1'b0 : free_adr_mask[143];
  assign free_adr_mask_next[143] = _2114_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:939" *) 1'b1 : _0221_;
  assign _0220_ = _2113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:936" *) 1'b0 : free_adr_mask[142];
  assign free_adr_mask_next[142] = _2112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:934" *) 1'b1 : _0220_;
  assign _0219_ = _2111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:931" *) 1'b0 : free_adr_mask[141];
  assign free_adr_mask_next[141] = _2110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:929" *) 1'b1 : _0219_;
  assign _0218_ = _2109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:926" *) 1'b0 : free_adr_mask[140];
  assign free_adr_mask_next[140] = _2108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:924" *) 1'b1 : _0218_;
  assign _0217_ = _2107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:921" *) 1'b0 : free_adr_mask[139];
  assign free_adr_mask_next[139] = _2106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:919" *) 1'b1 : _0217_;
  assign _0216_ = _2105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:916" *) 1'b0 : free_adr_mask[138];
  assign free_adr_mask_next[138] = _2104_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:914" *) 1'b1 : _0216_;
  assign _0215_ = _2103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:911" *) 1'b0 : free_adr_mask[137];
  assign free_adr_mask_next[137] = _2102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:909" *) 1'b1 : _0215_;
  assign _0214_ = _2101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:906" *) 1'b0 : free_adr_mask[136];
  assign free_adr_mask_next[136] = _2100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:904" *) 1'b1 : _0214_;
  assign _0213_ = _2099_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:901" *) 1'b0 : free_adr_mask[135];
  assign free_adr_mask_next[135] = _2098_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:899" *) 1'b1 : _0213_;
  assign _0212_ = _2097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:896" *) 1'b0 : free_adr_mask[134];
  assign free_adr_mask_next[134] = _2096_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:894" *) 1'b1 : _0212_;
  assign _0210_ = _2095_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:891" *) 1'b0 : free_adr_mask[133];
  assign free_adr_mask_next[133] = _2094_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:889" *) 1'b1 : _0210_;
  assign _0209_ = _2093_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:886" *) 1'b0 : free_adr_mask[132];
  assign free_adr_mask_next[132] = _2092_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:884" *) 1'b1 : _0209_;
  assign _0208_ = _2091_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:881" *) 1'b0 : free_adr_mask[131];
  assign free_adr_mask_next[131] = _2090_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:879" *) 1'b1 : _0208_;
  assign _0207_ = _2089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:876" *) 1'b0 : free_adr_mask[130];
  assign free_adr_mask_next[130] = _2088_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:874" *) 1'b1 : _0207_;
  assign _0206_ = _2087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:871" *) 1'b0 : free_adr_mask[129];
  assign free_adr_mask_next[129] = _2086_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:869" *) 1'b1 : _0206_;
  assign _0205_ = _2085_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:866" *) 1'b0 : free_adr_mask[128];
  assign free_adr_mask_next[128] = _2084_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:864" *) 1'b1 : _0205_;
  assign _0204_ = _2083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:861" *) 1'b0 : free_adr_mask[127];
  assign free_adr_mask_next[127] = _2082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:859" *) 1'b1 : _0204_;
  assign _0203_ = _2081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:856" *) 1'b0 : free_adr_mask[126];
  assign free_adr_mask_next[126] = _2080_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:854" *) 1'b1 : _0203_;
  assign _0202_ = _2079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:851" *) 1'b0 : free_adr_mask[125];
  assign free_adr_mask_next[125] = _2078_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:849" *) 1'b1 : _0202_;
  assign _0201_ = _2077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:846" *) 1'b0 : free_adr_mask[124];
  assign free_adr_mask_next[124] = _2076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:844" *) 1'b1 : _0201_;
  assign _0199_ = _2075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:841" *) 1'b0 : free_adr_mask[123];
  assign free_adr_mask_next[123] = _2074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:839" *) 1'b1 : _0199_;
  assign _0198_ = _2073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:836" *) 1'b0 : free_adr_mask[122];
  assign free_adr_mask_next[122] = _2072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:834" *) 1'b1 : _0198_;
  assign _0197_ = _2071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:831" *) 1'b0 : free_adr_mask[121];
  assign free_adr_mask_next[121] = _2070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:829" *) 1'b1 : _0197_;
  assign _0196_ = _2069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:826" *) 1'b0 : free_adr_mask[120];
  assign free_adr_mask_next[120] = _2068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:824" *) 1'b1 : _0196_;
  assign _0195_ = _2067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:821" *) 1'b0 : free_adr_mask[119];
  assign free_adr_mask_next[119] = _2066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:819" *) 1'b1 : _0195_;
  assign _0194_ = _2065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:816" *) 1'b0 : free_adr_mask[118];
  assign free_adr_mask_next[118] = _2064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:814" *) 1'b1 : _0194_;
  assign _0193_ = _2063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:811" *) 1'b0 : free_adr_mask[117];
  assign free_adr_mask_next[117] = _2062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:809" *) 1'b1 : _0193_;
  assign _0192_ = _2061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:806" *) 1'b0 : free_adr_mask[116];
  assign free_adr_mask_next[116] = _2060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:804" *) 1'b1 : _0192_;
  assign _0191_ = _2059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:801" *) 1'b0 : free_adr_mask[115];
  assign free_adr_mask_next[115] = _2058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:799" *) 1'b1 : _0191_;
  assign _0190_ = _2057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:796" *) 1'b0 : free_adr_mask[114];
  assign free_adr_mask_next[114] = _2056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:794" *) 1'b1 : _0190_;
  assign _0188_ = _2055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:791" *) 1'b0 : free_adr_mask[113];
  assign free_adr_mask_next[113] = _2054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:789" *) 1'b1 : _0188_;
  assign _0187_ = _2053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:786" *) 1'b0 : free_adr_mask[112];
  assign free_adr_mask_next[112] = _2052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:784" *) 1'b1 : _0187_;
  assign _0186_ = _2051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:781" *) 1'b0 : free_adr_mask[111];
  assign free_adr_mask_next[111] = _2050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:779" *) 1'b1 : _0186_;
  assign _0185_ = _2049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:776" *) 1'b0 : free_adr_mask[110];
  assign free_adr_mask_next[110] = _2048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:774" *) 1'b1 : _0185_;
  assign _0184_ = _2047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:771" *) 1'b0 : free_adr_mask[109];
  assign free_adr_mask_next[109] = _2046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:769" *) 1'b1 : _0184_;
  assign _0183_ = _2045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:766" *) 1'b0 : free_adr_mask[108];
  assign free_adr_mask_next[108] = _2044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:764" *) 1'b1 : _0183_;
  assign _0182_ = _2043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:761" *) 1'b0 : free_adr_mask[107];
  assign free_adr_mask_next[107] = _2042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:759" *) 1'b1 : _0182_;
  assign _0181_ = _2041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:756" *) 1'b0 : free_adr_mask[106];
  assign free_adr_mask_next[106] = _2040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:754" *) 1'b1 : _0181_;
  assign _0180_ = _2039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:751" *) 1'b0 : free_adr_mask[105];
  assign free_adr_mask_next[105] = _2038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:749" *) 1'b1 : _0180_;
  assign _0179_ = _2037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:746" *) 1'b0 : free_adr_mask[104];
  assign free_adr_mask_next[104] = _2036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:744" *) 1'b1 : _0179_;
  assign _0177_ = _2035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:741" *) 1'b0 : free_adr_mask[103];
  assign free_adr_mask_next[103] = _2034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:739" *) 1'b1 : _0177_;
  assign _0176_ = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:736" *) 1'b0 : free_adr_mask[102];
  assign free_adr_mask_next[102] = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:734" *) 1'b1 : _0176_;
  assign _0175_ = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:731" *) 1'b0 : free_adr_mask[101];
  assign free_adr_mask_next[101] = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:729" *) 1'b1 : _0175_;
  assign _0174_ = _2029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:726" *) 1'b0 : free_adr_mask[100];
  assign free_adr_mask_next[100] = _2028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:724" *) 1'b1 : _0174_;
  assign _0173_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:721" *) 1'b0 : free_adr_mask[99];
  assign free_adr_mask_next[99] = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:719" *) 1'b1 : _0173_;
  assign _0172_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:716" *) 1'b0 : free_adr_mask[98];
  assign free_adr_mask_next[98] = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:714" *) 1'b1 : _0172_;
  assign _0171_ = _2023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:711" *) 1'b0 : free_adr_mask[97];
  assign free_adr_mask_next[97] = _2022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:709" *) 1'b1 : _0171_;
  assign _0170_ = _2021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:706" *) 1'b0 : free_adr_mask[96];
  assign free_adr_mask_next[96] = _2020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:704" *) 1'b1 : _0170_;
  assign _0169_ = _2019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:701" *) 1'b0 : free_adr_mask[95];
  assign free_adr_mask_next[95] = _2018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:699" *) 1'b1 : _0169_;
  assign _0168_ = _2017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:696" *) 1'b0 : free_adr_mask[94];
  assign free_adr_mask_next[94] = _2016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:694" *) 1'b1 : _0168_;
  assign _0166_ = _2015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:691" *) 1'b0 : free_adr_mask[93];
  assign free_adr_mask_next[93] = _2014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:689" *) 1'b1 : _0166_;
  assign _0165_ = _2013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:686" *) 1'b0 : free_adr_mask[92];
  assign free_adr_mask_next[92] = _2012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:684" *) 1'b1 : _0165_;
  assign _0164_ = _2011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:681" *) 1'b0 : free_adr_mask[91];
  assign free_adr_mask_next[91] = _2010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:679" *) 1'b1 : _0164_;
  assign _0163_ = _2009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:676" *) 1'b0 : free_adr_mask[90];
  assign free_adr_mask_next[90] = _2008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:674" *) 1'b1 : _0163_;
  assign _0162_ = _2007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:671" *) 1'b0 : free_adr_mask[89];
  assign free_adr_mask_next[89] = _2006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:669" *) 1'b1 : _0162_;
  assign _0161_ = _2005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:666" *) 1'b0 : free_adr_mask[88];
  assign free_adr_mask_next[88] = _2004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:664" *) 1'b1 : _0161_;
  assign _0160_ = _2003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:661" *) 1'b0 : free_adr_mask[87];
  assign free_adr_mask_next[87] = _2002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:659" *) 1'b1 : _0160_;
  assign _0159_ = _2001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:656" *) 1'b0 : free_adr_mask[86];
  assign free_adr_mask_next[86] = _2000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:654" *) 1'b1 : _0159_;
  assign _0158_ = _1999_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:651" *) 1'b0 : free_adr_mask[85];
  assign free_adr_mask_next[85] = _1998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:649" *) 1'b1 : _0158_;
  assign _0157_ = _1997_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:646" *) 1'b0 : free_adr_mask[84];
  assign free_adr_mask_next[84] = _1996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:644" *) 1'b1 : _0157_;
  assign _0155_ = _1995_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:641" *) 1'b0 : free_adr_mask[83];
  assign free_adr_mask_next[83] = _1994_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:639" *) 1'b1 : _0155_;
  assign _0154_ = _1993_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:636" *) 1'b0 : free_adr_mask[82];
  assign free_adr_mask_next[82] = _1992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:634" *) 1'b1 : _0154_;
  assign _0153_ = _1991_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:631" *) 1'b0 : free_adr_mask[81];
  assign free_adr_mask_next[81] = _1990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:629" *) 1'b1 : _0153_;
  assign _0152_ = _1989_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:626" *) 1'b0 : free_adr_mask[80];
  assign free_adr_mask_next[80] = _1988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:624" *) 1'b1 : _0152_;
  assign _0151_ = _1987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:621" *) 1'b0 : free_adr_mask[79];
  assign free_adr_mask_next[79] = _1986_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:619" *) 1'b1 : _0151_;
  assign _0150_ = _1985_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:616" *) 1'b0 : free_adr_mask[78];
  assign free_adr_mask_next[78] = _1984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:614" *) 1'b1 : _0150_;
  assign _0149_ = _1983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:611" *) 1'b0 : free_adr_mask[77];
  assign free_adr_mask_next[77] = _1982_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:609" *) 1'b1 : _0149_;
  assign _0148_ = _1981_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:606" *) 1'b0 : free_adr_mask[76];
  assign free_adr_mask_next[76] = _1980_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:604" *) 1'b1 : _0148_;
  assign _0147_ = _1979_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:601" *) 1'b0 : free_adr_mask[75];
  assign free_adr_mask_next[75] = _1978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:599" *) 1'b1 : _0147_;
  assign _0146_ = _1977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:596" *) 1'b0 : free_adr_mask[74];
  assign free_adr_mask_next[74] = _1976_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:594" *) 1'b1 : _0146_;
  assign _0144_ = _1975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:591" *) 1'b0 : free_adr_mask[73];
  assign free_adr_mask_next[73] = _1974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:589" *) 1'b1 : _0144_;
  assign _0143_ = _1973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:586" *) 1'b0 : free_adr_mask[72];
  assign free_adr_mask_next[72] = _1972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:584" *) 1'b1 : _0143_;
  assign _0142_ = _1971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:581" *) 1'b0 : free_adr_mask[71];
  assign free_adr_mask_next[71] = _1970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:579" *) 1'b1 : _0142_;
  assign _0141_ = _1969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:576" *) 1'b0 : free_adr_mask[70];
  assign free_adr_mask_next[70] = _1968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:574" *) 1'b1 : _0141_;
  assign _0140_ = _1967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:571" *) 1'b0 : free_adr_mask[69];
  assign free_adr_mask_next[69] = _1966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:569" *) 1'b1 : _0140_;
  assign _0139_ = _1965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:566" *) 1'b0 : free_adr_mask[68];
  assign free_adr_mask_next[68] = _1964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:564" *) 1'b1 : _0139_;
  assign _0138_ = _1963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:561" *) 1'b0 : free_adr_mask[67];
  assign free_adr_mask_next[67] = _1962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:559" *) 1'b1 : _0138_;
  assign _0137_ = _1961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:556" *) 1'b0 : free_adr_mask[66];
  assign free_adr_mask_next[66] = _1960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:554" *) 1'b1 : _0137_;
  assign _0136_ = _1959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:551" *) 1'b0 : free_adr_mask[65];
  assign free_adr_mask_next[65] = _1958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:549" *) 1'b1 : _0136_;
  assign _0135_ = _1957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:546" *) 1'b0 : free_adr_mask[64];
  assign free_adr_mask_next[64] = _1956_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:544" *) 1'b1 : _0135_;
  assign _0133_ = _1955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:541" *) 1'b0 : free_adr_mask[63];
  assign free_adr_mask_next[63] = _1954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:539" *) 1'b1 : _0133_;
  assign _0132_ = _1953_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:536" *) 1'b0 : free_adr_mask[62];
  assign free_adr_mask_next[62] = _1952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:534" *) 1'b1 : _0132_;
  assign _0131_ = _1951_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:531" *) 1'b0 : free_adr_mask[61];
  assign free_adr_mask_next[61] = _1950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:529" *) 1'b1 : _0131_;
  assign _0130_ = _1949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:526" *) 1'b0 : free_adr_mask[60];
  assign free_adr_mask_next[60] = _1948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:524" *) 1'b1 : _0130_;
  assign _0129_ = _1947_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:521" *) 1'b0 : free_adr_mask[59];
  assign free_adr_mask_next[59] = _1946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:519" *) 1'b1 : _0129_;
  assign _0128_ = _1945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:516" *) 1'b0 : free_adr_mask[58];
  assign free_adr_mask_next[58] = _1944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:514" *) 1'b1 : _0128_;
  assign _0127_ = _1943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:511" *) 1'b0 : free_adr_mask[57];
  assign free_adr_mask_next[57] = _1942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:509" *) 1'b1 : _0127_;
  assign _0126_ = _1941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:506" *) 1'b0 : free_adr_mask[56];
  assign free_adr_mask_next[56] = _1940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:504" *) 1'b1 : _0126_;
  assign _0125_ = _1939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:501" *) 1'b0 : free_adr_mask[55];
  assign free_adr_mask_next[55] = _1938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:499" *) 1'b1 : _0125_;
  assign _0124_ = _1937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:496" *) 1'b0 : free_adr_mask[54];
  assign free_adr_mask_next[54] = _1936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:494" *) 1'b1 : _0124_;
  assign _0122_ = _1935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:491" *) 1'b0 : free_adr_mask[53];
  assign free_adr_mask_next[53] = _1934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:489" *) 1'b1 : _0122_;
  assign _0121_ = _1933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:486" *) 1'b0 : free_adr_mask[52];
  assign free_adr_mask_next[52] = _1932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:484" *) 1'b1 : _0121_;
  assign _0120_ = _1931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:481" *) 1'b0 : free_adr_mask[51];
  assign free_adr_mask_next[51] = _1930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:479" *) 1'b1 : _0120_;
  assign _0119_ = _1929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:476" *) 1'b0 : free_adr_mask[50];
  assign free_adr_mask_next[50] = _1928_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:474" *) 1'b1 : _0119_;
  assign _0118_ = _1927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:471" *) 1'b0 : free_adr_mask[49];
  assign free_adr_mask_next[49] = _1926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:469" *) 1'b1 : _0118_;
  assign _0372_ = _1925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:466" *) 1'b0 : free_adr_mask[48];
  assign free_adr_mask_next[48] = _1924_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:464" *) 1'b1 : _0372_;
  assign _0371_ = _1923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:461" *) 1'b0 : free_adr_mask[47];
  assign free_adr_mask_next[47] = _1922_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:459" *) 1'b1 : _0371_;
  assign _0370_ = _1921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:456" *) 1'b0 : free_adr_mask[46];
  assign free_adr_mask_next[46] = _1920_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:454" *) 1'b1 : _0370_;
  assign _0369_ = _1919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:451" *) 1'b0 : free_adr_mask[45];
  assign free_adr_mask_next[45] = _1918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:449" *) 1'b1 : _0369_;
  assign _0368_ = _1917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:446" *) 1'b0 : free_adr_mask[44];
  assign free_adr_mask_next[44] = _1916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:444" *) 1'b1 : _0368_;
  assign _0366_ = _1915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:441" *) 1'b0 : free_adr_mask[43];
  assign free_adr_mask_next[43] = _1914_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:439" *) 1'b1 : _0366_;
  assign _0365_ = _1913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:436" *) 1'b0 : free_adr_mask[42];
  assign free_adr_mask_next[42] = _1912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:434" *) 1'b1 : _0365_;
  assign _0364_ = _1911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:431" *) 1'b0 : free_adr_mask[41];
  assign free_adr_mask_next[41] = _1910_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:429" *) 1'b1 : _0364_;
  assign _0363_ = _1909_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:426" *) 1'b0 : free_adr_mask[40];
  assign free_adr_mask_next[40] = _1908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:424" *) 1'b1 : _0363_;
  assign _0362_ = _1907_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:421" *) 1'b0 : free_adr_mask[39];
  assign free_adr_mask_next[39] = _1906_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:419" *) 1'b1 : _0362_;
  assign _0361_ = _1905_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:416" *) 1'b0 : free_adr_mask[38];
  assign free_adr_mask_next[38] = _1904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:414" *) 1'b1 : _0361_;
  assign _0360_ = _1903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:411" *) 1'b0 : free_adr_mask[37];
  assign free_adr_mask_next[37] = _1902_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:409" *) 1'b1 : _0360_;
  assign _0359_ = _1901_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:406" *) 1'b0 : free_adr_mask[36];
  assign free_adr_mask_next[36] = _1900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:404" *) 1'b1 : _0359_;
  assign _0358_ = _1899_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:401" *) 1'b0 : free_adr_mask[35];
  assign free_adr_mask_next[35] = _1898_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:399" *) 1'b1 : _0358_;
  assign _0357_ = _1897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:396" *) 1'b0 : free_adr_mask[34];
  assign free_adr_mask_next[34] = _1896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:394" *) 1'b1 : _0357_;
  assign _0355_ = _1895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:391" *) 1'b0 : free_adr_mask[33];
  assign free_adr_mask_next[33] = _1894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:389" *) 1'b1 : _0355_;
  assign _0354_ = _1893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:386" *) 1'b0 : free_adr_mask[32];
  assign free_adr_mask_next[32] = _1892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:384" *) 1'b1 : _0354_;
  assign _0353_ = _1891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:381" *) 1'b0 : free_adr_mask[31];
  assign free_adr_mask_next[31] = _1890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:379" *) 1'b1 : _0353_;
  assign _0352_ = _1889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:376" *) 1'b0 : free_adr_mask[30];
  assign free_adr_mask_next[30] = _1888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:374" *) 1'b1 : _0352_;
  assign _0351_ = _1887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:371" *) 1'b0 : free_adr_mask[29];
  assign free_adr_mask_next[29] = _1886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:369" *) 1'b1 : _0351_;
  assign _0350_ = _1885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:366" *) 1'b0 : free_adr_mask[28];
  assign free_adr_mask_next[28] = _1884_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:364" *) 1'b1 : _0350_;
  assign _0349_ = _1875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:361" *) 1'b0 : free_adr_mask[27];
  assign free_adr_mask_next[27] = _1792_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:359" *) 1'b1 : _0349_;
  assign _0348_ = _1674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:356" *) 1'b0 : free_adr_mask[26];
  assign free_adr_mask_next[26] = _1590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:354" *) 1'b1 : _0348_;
  assign _0347_ = _1474_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:351" *) 1'b0 : free_adr_mask[25];
  assign free_adr_mask_next[25] = _1467_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:349" *) 1'b1 : _0347_;
  assign _0345_ = _1462_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:346" *) 1'b0 : free_adr_mask[24];
  assign free_adr_mask_next[24] = _1455_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:344" *) 1'b1 : _0345_;
  assign _0333_ = _1450_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:341" *) 1'b0 : free_adr_mask[23];
  assign free_adr_mask_next[23] = _1442_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:339" *) 1'b1 : _0333_;
  assign _0322_ = _1435_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:336" *) 1'b0 : free_adr_mask[22];
  assign free_adr_mask_next[22] = _1431_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:334" *) 1'b1 : _0322_;
  assign _0311_ = _1426_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:331" *) 1'b0 : free_adr_mask[21];
  assign free_adr_mask_next[21] = _1418_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:329" *) 1'b1 : _0311_;
  assign _0300_ = _1411_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:326" *) 1'b0 : free_adr_mask[20];
  assign free_adr_mask_next[20] = _1403_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:324" *) 1'b1 : _0300_;
  assign _0289_ = _1402_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:321" *) 1'b0 : free_adr_mask[19];
  assign free_adr_mask_next[19] = _1394_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:319" *) 1'b1 : _0289_;
  assign _0278_ = _1387_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:316" *) 1'b0 : free_adr_mask[18];
  assign free_adr_mask_next[18] = _1379_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:314" *) 1'b1 : _0278_;
  assign _0267_ = _1378_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:311" *) 1'b0 : free_adr_mask[17];
  assign free_adr_mask_next[17] = _1368_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:309" *) 1'b1 : _0267_;
  assign _0256_ = _1360_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:306" *) 1'b0 : free_adr_mask[16];
  assign free_adr_mask_next[16] = _1355_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:304" *) 1'b1 : _0256_;
  assign _0245_ = _1348_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:301" *) 1'b0 : free_adr_mask[15];
  assign free_adr_mask_next[15] = _1343_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:299" *) 1'b1 : _0245_;
  assign _0234_ = _1336_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:296" *) 1'b0 : free_adr_mask[14];
  assign free_adr_mask_next[14] = _1331_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:294" *) 1'b1 : _0234_;
  assign _0222_ = _1323_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:291" *) 1'b0 : free_adr_mask[13];
  assign free_adr_mask_next[13] = _1319_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:289" *) 1'b1 : _0222_;
  assign _0211_ = _1312_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:286" *) 1'b0 : free_adr_mask[12];
  assign free_adr_mask_next[12] = _1307_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:284" *) 1'b1 : _0211_;
  assign _0200_ = _1299_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:281" *) 1'b0 : free_adr_mask[11];
  assign free_adr_mask_next[11] = _1295_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:279" *) 1'b1 : _0200_;
  assign _0189_ = _1284_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:276" *) 1'b0 : free_adr_mask[10];
  assign free_adr_mask_next[10] = _1283_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:274" *) 1'b1 : _0189_;
  assign _0178_ = _1275_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:271" *) 1'b0 : free_adr_mask[9];
  assign free_adr_mask_next[9] = _1271_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:269" *) 1'b1 : _0178_;
  assign _0167_ = _1260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:266" *) 1'b0 : free_adr_mask[8];
  assign free_adr_mask_next[8] = _1259_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:264" *) 1'b1 : _0167_;
  assign _0156_ = _1249_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:261" *) 1'b0 : free_adr_mask[7];
  assign free_adr_mask_next[7] = _1244_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:259" *) 1'b1 : _0156_;
  assign _0145_ = _1236_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:256" *) 1'b0 : free_adr_mask[6];
  assign free_adr_mask_next[6] = _1235_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:254" *) 1'b1 : _0145_;
  assign _0134_ = _1234_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:251" *) 1'b0 : free_adr_mask[5];
  assign free_adr_mask_next[5] = _1223_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:249" *) 1'b1 : _0134_;
  assign _0123_ = _1205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:246" *) 1'b0 : free_adr_mask[4];
  assign free_adr_mask_next[4] = _1201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:244" *) 1'b1 : _0123_;
  assign _0367_ = _1197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:241" *) 1'b0 : free_adr_mask[3];
  assign free_adr_mask_next[3] = _1190_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:239" *) 1'b1 : _0367_;
  assign _0356_ = _1183_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:236" *) 1'b0 : free_adr_mask[2];
  assign free_adr_mask_next[2] = _1179_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:234" *) 1'b1 : _0356_;
  assign _0339_ = _1172_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:231" *) 1'b0 : free_adr_mask[1];
  assign free_adr_mask_next[1] = _1168_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:229" *) 1'b1 : _0339_;
  assign _0228_ = _1164_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:226" *) 1'b0 : free_adr_mask[0];
  assign free_adr_mask_next[0] = _1163_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:224" *) 1'b1 : _0228_;
  assign _0033_ = _2231_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:211" *) free_adr_mask_next : free_adr_mask;
  assign _0032_ = _2529_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:162" *) wr_count_next : cq_wr_count;
  assign cq_rd_take = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3510" *) { cq_rd_take_elig[0], cq_rd_take_elig[1], cq_rd_take_elig[2], cq_rd_take_elig[3], cq_rd_take_elig[4], cq_rd_take_elig[5], cq_rd_take_elig[6], cq_rd_take_elig[7], cq_rd_take_elig[8], cq_rd_take_elig[9] };
  assign cq_rd_take_thread_id[0] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3611" *) { cq_rd_take_thread_id_is_1[0], cq_rd_take_thread_id_is_1[1], cq_rd_take_thread_id_is_1[2], cq_rd_take_thread_id_is_1[3], cq_rd_take_thread_id_is_1[4], cq_rd_take_thread_id_is_1[5], cq_rd_take_thread_id_is_1[6], cq_rd_take_thread_id_is_1[7], cq_rd_take_thread_id_is_1[8], cq_rd_take_thread_id_is_1[9], cq_rd_take_thread_id_is_3[0], cq_rd_take_thread_id_is_3[1], cq_rd_take_thread_id_is_3[2], cq_rd_take_thread_id_is_3[3], cq_rd_take_thread_id_is_3[4], cq_rd_take_thread_id_is_3[5], cq_rd_take_thread_id_is_3[6], cq_rd_take_thread_id_is_3[7], cq_rd_take_thread_id_is_3[8], cq_rd_take_thread_id_is_3[9], cq_rd_take_thread_id_is_5[0], cq_rd_take_thread_id_is_5[1], cq_rd_take_thread_id_is_5[2], cq_rd_take_thread_id_is_5[3], cq_rd_take_thread_id_is_5[4], cq_rd_take_thread_id_is_5[5], cq_rd_take_thread_id_is_5[6], cq_rd_take_thread_id_is_5[7], cq_rd_take_thread_id_is_5[8], cq_rd_take_thread_id_is_5[9], cq_rd_take_thread_id_is_7[0], cq_rd_take_thread_id_is_7[1], cq_rd_take_thread_id_is_7[2], cq_rd_take_thread_id_is_7[3], cq_rd_take_thread_id_is_7[4], cq_rd_take_thread_id_is_7[5], cq_rd_take_thread_id_is_7[6], cq_rd_take_thread_id_is_7[7], cq_rd_take_thread_id_is_7[8], cq_rd_take_thread_id_is_7[9], cq_rd_take_thread_id_is_9[0], cq_rd_take_thread_id_is_9[1], cq_rd_take_thread_id_is_9[2], cq_rd_take_thread_id_is_9[3], cq_rd_take_thread_id_is_9[4], cq_rd_take_thread_id_is_9[5], cq_rd_take_thread_id_is_9[6], cq_rd_take_thread_id_is_9[7], cq_rd_take_thread_id_is_9[8], cq_rd_take_thread_id_is_9[9] };
  assign cq_rd_take_thread_id[1] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3612" *) { cq_rd_take_thread_id_is_2[0], cq_rd_take_thread_id_is_2[1], cq_rd_take_thread_id_is_2[2], cq_rd_take_thread_id_is_2[3], cq_rd_take_thread_id_is_2[4], cq_rd_take_thread_id_is_2[5], cq_rd_take_thread_id_is_2[6], cq_rd_take_thread_id_is_2[7], cq_rd_take_thread_id_is_2[8], cq_rd_take_thread_id_is_2[9], cq_rd_take_thread_id_is_3[0], cq_rd_take_thread_id_is_3[1], cq_rd_take_thread_id_is_3[2], cq_rd_take_thread_id_is_3[3], cq_rd_take_thread_id_is_3[4], cq_rd_take_thread_id_is_3[5], cq_rd_take_thread_id_is_3[6], cq_rd_take_thread_id_is_3[7], cq_rd_take_thread_id_is_3[8], cq_rd_take_thread_id_is_3[9], cq_rd_take_thread_id_is_6[0], cq_rd_take_thread_id_is_6[1], cq_rd_take_thread_id_is_6[2], cq_rd_take_thread_id_is_6[3], cq_rd_take_thread_id_is_6[4], cq_rd_take_thread_id_is_6[5], cq_rd_take_thread_id_is_6[6], cq_rd_take_thread_id_is_6[7], cq_rd_take_thread_id_is_6[8], cq_rd_take_thread_id_is_6[9], cq_rd_take_thread_id_is_7[0], cq_rd_take_thread_id_is_7[1], cq_rd_take_thread_id_is_7[2], cq_rd_take_thread_id_is_7[3], cq_rd_take_thread_id_is_7[4], cq_rd_take_thread_id_is_7[5], cq_rd_take_thread_id_is_7[6], cq_rd_take_thread_id_is_7[7], cq_rd_take_thread_id_is_7[8], cq_rd_take_thread_id_is_7[9] };
  assign cq_rd_take_thread_id[2] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3613" *) { cq_rd_take_thread_id_is_4[0], cq_rd_take_thread_id_is_4[1], cq_rd_take_thread_id_is_4[2], cq_rd_take_thread_id_is_4[3], cq_rd_take_thread_id_is_4[4], cq_rd_take_thread_id_is_4[5], cq_rd_take_thread_id_is_4[6], cq_rd_take_thread_id_is_4[7], cq_rd_take_thread_id_is_4[8], cq_rd_take_thread_id_is_4[9], cq_rd_take_thread_id_is_5[0], cq_rd_take_thread_id_is_5[1], cq_rd_take_thread_id_is_5[2], cq_rd_take_thread_id_is_5[3], cq_rd_take_thread_id_is_5[4], cq_rd_take_thread_id_is_5[5], cq_rd_take_thread_id_is_5[6], cq_rd_take_thread_id_is_5[7], cq_rd_take_thread_id_is_5[8], cq_rd_take_thread_id_is_5[9], cq_rd_take_thread_id_is_6[0], cq_rd_take_thread_id_is_6[1], cq_rd_take_thread_id_is_6[2], cq_rd_take_thread_id_is_6[3], cq_rd_take_thread_id_is_6[4], cq_rd_take_thread_id_is_6[5], cq_rd_take_thread_id_is_6[6], cq_rd_take_thread_id_is_6[7], cq_rd_take_thread_id_is_6[8], cq_rd_take_thread_id_is_6[9], cq_rd_take_thread_id_is_7[0], cq_rd_take_thread_id_is_7[1], cq_rd_take_thread_id_is_7[2], cq_rd_take_thread_id_is_7[3], cq_rd_take_thread_id_is_7[4], cq_rd_take_thread_id_is_7[5], cq_rd_take_thread_id_is_7[6], cq_rd_take_thread_id_is_7[7], cq_rd_take_thread_id_is_7[8], cq_rd_take_thread_id_is_7[9] };
  assign cq_rd_take_thread_id[3] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3614" *) { cq_rd_take_thread_id_is_8[0], cq_rd_take_thread_id_is_8[1], cq_rd_take_thread_id_is_8[2], cq_rd_take_thread_id_is_8[3], cq_rd_take_thread_id_is_8[4], cq_rd_take_thread_id_is_8[5], cq_rd_take_thread_id_is_8[6], cq_rd_take_thread_id_is_8[7], cq_rd_take_thread_id_is_8[8], cq_rd_take_thread_id_is_8[9], cq_rd_take_thread_id_is_9[0], cq_rd_take_thread_id_is_9[1], cq_rd_take_thread_id_is_9[2], cq_rd_take_thread_id_is_9[3], cq_rd_take_thread_id_is_9[4], cq_rd_take_thread_id_is_9[5], cq_rd_take_thread_id_is_9[6], cq_rd_take_thread_id_is_9[7], cq_rd_take_thread_id_is_9[8], cq_rd_take_thread_id_is_9[9] };
  assign _2530_ = cq_wr_count - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:126" *) 1'b1;
  assign _2531_ = cq_rd_count0 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2115" *) 1'b1;
  assign _2532_ = cq_rd_count1 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2118" *) 1'b1;
  assign _2533_ = cq_rd_count2 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2121" *) 1'b1;
  assign _2534_ = cq_rd_count3 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2124" *) 1'b1;
  assign _2535_ = cq_rd_count4 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2127" *) 1'b1;
  assign _2536_ = cq_rd_count5 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2130" *) 1'b1;
  assign _2537_ = cq_rd_count6 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2133" *) 1'b1;
  assign _2538_ = cq_rd_count7 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2136" *) 1'b1;
  assign _2539_ = cq_rd_count8 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2139" *) 1'b1;
  assign _2540_ = cq_rd_count9 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2142" *) 1'b1;
  assign cq_rd0_credits_w_take_next = cq_rd0_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2619" *) 1'b1;
  assign cq_rd1_credits_w_take_next = cq_rd1_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2715" *) 1'b1;
  assign cq_rd2_credits_w_take_next = cq_rd2_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2811" *) 1'b1;
  assign cq_rd3_credits_w_take_next = cq_rd3_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2907" *) 1'b1;
  assign cq_rd4_credits_w_take_next = cq_rd4_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3003" *) 1'b1;
  assign cq_rd5_credits_w_take_next = cq_rd5_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3099" *) 1'b1;
  assign cq_rd6_credits_w_take_next = cq_rd6_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3195" *) 1'b1;
  assign cq_rd7_credits_w_take_next = cq_rd7_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3291" *) 1'b1;
  assign cq_rd8_credits_w_take_next = cq_rd8_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3387" *) 1'b1;
  assign cq_rd9_credits_w_take_next = cq_rd9_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3483" *) 1'b1;
  assign wr_count_next_wr_popping = rd_pushing ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:126" *) cq_wr_count : _2530_;
  assign wr_count_next_no_wr_popping = rd_pushing ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:127" *) _0373_ : cq_wr_count;
  assign wr_count_next = rd_take_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:129" *) wr_count_next_wr_popping : wr_count_next_no_wr_popping;
  assign cq_wr_busy_next = rd_take_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:132" *) 1'b0 : wr_count_next_no_wr_popping_is_256;
  assign index_l1_0[0] = flag_l0_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1875" *) index_l0_0 : index_l0_1;
  assign index_l1_1[0] = flag_l0_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1876" *) index_l0_2 : index_l0_3;
  assign index_l1_2[0] = flag_l0_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1877" *) index_l0_4 : index_l0_5;
  assign index_l1_3[0] = flag_l0_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1878" *) index_l0_6 : index_l0_7;
  assign index_l1_4[0] = flag_l0_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1879" *) index_l0_8 : index_l0_9;
  assign index_l1_5[0] = flag_l0_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1880" *) index_l0_10 : index_l0_11;
  assign index_l1_6[0] = flag_l0_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1881" *) index_l0_12 : index_l0_13;
  assign index_l1_7[0] = flag_l0_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1882" *) index_l0_14 : index_l0_15;
  assign index_l1_8[0] = flag_l0_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1883" *) index_l0_16 : index_l0_17;
  assign index_l1_9[0] = flag_l0_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1884" *) index_l0_18 : index_l0_19;
  assign index_l1_10[0] = flag_l0_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1885" *) index_l0_20 : index_l0_21;
  assign index_l1_11[0] = flag_l0_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1886" *) index_l0_22 : index_l0_23;
  assign index_l1_12[0] = flag_l0_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1887" *) index_l0_24 : index_l0_25;
  assign index_l1_13[0] = flag_l0_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1888" *) index_l0_26 : index_l0_27;
  assign index_l1_14[0] = flag_l0_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1889" *) index_l0_28 : index_l0_29;
  assign index_l1_15[0] = flag_l0_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1890" *) index_l0_30 : index_l0_31;
  assign index_l1_16[0] = flag_l0_32 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1891" *) index_l0_32 : index_l0_33;
  assign index_l1_17[0] = flag_l0_34 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1892" *) index_l0_34 : index_l0_35;
  assign index_l1_18[0] = flag_l0_36 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1893" *) index_l0_36 : index_l0_37;
  assign index_l1_19[0] = flag_l0_38 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1894" *) index_l0_38 : index_l0_39;
  assign index_l1_20[0] = flag_l0_40 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1895" *) index_l0_40 : index_l0_41;
  assign index_l1_21[0] = flag_l0_42 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1896" *) index_l0_42 : index_l0_43;
  assign index_l1_22[0] = flag_l0_44 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1897" *) index_l0_44 : index_l0_45;
  assign index_l1_23[0] = flag_l0_46 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1898" *) index_l0_46 : index_l0_47;
  assign index_l1_24[0] = flag_l0_48 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1899" *) index_l0_48 : index_l0_49;
  assign index_l1_25[0] = flag_l0_50 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1900" *) index_l0_50 : index_l0_51;
  assign index_l1_26[0] = flag_l0_52 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1901" *) index_l0_52 : index_l0_53;
  assign index_l1_27[0] = flag_l0_54 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1902" *) index_l0_54 : index_l0_55;
  assign index_l1_28[0] = flag_l0_56 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1903" *) index_l0_56 : index_l0_57;
  assign index_l1_29[0] = flag_l0_58 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1904" *) index_l0_58 : index_l0_59;
  assign index_l1_30[0] = flag_l0_60 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1905" *) index_l0_60 : index_l0_61;
  assign index_l1_31[0] = flag_l0_62 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1906" *) index_l0_62 : index_l0_63;
  assign index_l1_32[0] = flag_l0_64 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1907" *) index_l0_64 : index_l0_65;
  assign index_l1_33[0] = flag_l0_66 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1908" *) index_l0_66 : index_l0_67;
  assign index_l1_34[0] = flag_l0_68 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1909" *) index_l0_68 : index_l0_69;
  assign index_l1_35[0] = flag_l0_70 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1910" *) index_l0_70 : index_l0_71;
  assign index_l1_36[0] = flag_l0_72 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1911" *) index_l0_72 : index_l0_73;
  assign index_l1_37[0] = flag_l0_74 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1912" *) index_l0_74 : index_l0_75;
  assign index_l1_38[0] = flag_l0_76 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1913" *) index_l0_76 : index_l0_77;
  assign index_l1_39[0] = flag_l0_78 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1914" *) index_l0_78 : index_l0_79;
  assign index_l1_40[0] = flag_l0_80 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1915" *) index_l0_80 : index_l0_81;
  assign index_l1_41[0] = flag_l0_82 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1916" *) index_l0_82 : index_l0_83;
  assign index_l1_42[0] = flag_l0_84 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1917" *) index_l0_84 : index_l0_85;
  assign index_l1_43[0] = flag_l0_86 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1918" *) index_l0_86 : index_l0_87;
  assign index_l1_44[0] = flag_l0_88 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1919" *) index_l0_88 : index_l0_89;
  assign index_l1_45[0] = flag_l0_90 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1920" *) index_l0_90 : index_l0_91;
  assign index_l1_46[0] = flag_l0_92 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1921" *) index_l0_92 : index_l0_93;
  assign index_l1_47[0] = flag_l0_94 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1922" *) index_l0_94 : index_l0_95;
  assign index_l1_48[0] = flag_l0_96 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1923" *) index_l0_96 : index_l0_97;
  assign index_l1_49[0] = flag_l0_98 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1924" *) index_l0_98 : index_l0_99;
  assign index_l1_50[0] = flag_l0_100 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1925" *) index_l0_100 : index_l0_101;
  assign index_l1_51[0] = flag_l0_102 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1926" *) index_l0_102 : index_l0_103;
  assign index_l1_52[0] = flag_l0_104 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1927" *) index_l0_104 : index_l0_105;
  assign index_l1_53[0] = flag_l0_106 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1928" *) index_l0_106 : index_l0_107;
  assign index_l1_54[0] = flag_l0_108 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1929" *) index_l0_108 : index_l0_109;
  assign index_l1_55[0] = flag_l0_110 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1930" *) index_l0_110 : index_l0_111;
  assign index_l1_56[0] = flag_l0_112 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1931" *) index_l0_112 : index_l0_113;
  assign index_l1_57[0] = flag_l0_114 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1932" *) index_l0_114 : index_l0_115;
  assign index_l1_58[0] = flag_l0_116 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1933" *) index_l0_116 : index_l0_117;
  assign index_l1_59[0] = flag_l0_118 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1934" *) index_l0_118 : index_l0_119;
  assign index_l1_60[0] = flag_l0_120 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1935" *) index_l0_120 : index_l0_121;
  assign index_l1_61[0] = flag_l0_122 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1936" *) index_l0_122 : index_l0_123;
  assign index_l1_62[0] = flag_l0_124 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1937" *) index_l0_124 : index_l0_125;
  assign index_l1_63[0] = flag_l0_126 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1938" *) index_l0_126 : index_l0_127;
  assign index_l2_0[1:0] = flag_l1_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1939" *) index_l1_0 : index_l1_1;
  assign index_l2_1[1:0] = flag_l1_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1940" *) index_l1_2 : index_l1_3;
  assign index_l2_2[1:0] = flag_l1_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1941" *) index_l1_4 : index_l1_5;
  assign index_l2_3[1:0] = flag_l1_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1942" *) index_l1_6 : index_l1_7;
  assign index_l2_4[1:0] = flag_l1_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1943" *) index_l1_8 : index_l1_9;
  assign index_l2_5[1:0] = flag_l1_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1944" *) index_l1_10 : index_l1_11;
  assign index_l2_6[1:0] = flag_l1_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1945" *) index_l1_12 : index_l1_13;
  assign index_l2_7[1:0] = flag_l1_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1946" *) index_l1_14 : index_l1_15;
  assign index_l2_8[1:0] = flag_l1_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1947" *) index_l1_16 : index_l1_17;
  assign index_l2_9[1:0] = flag_l1_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1948" *) index_l1_18 : index_l1_19;
  assign index_l2_10[1:0] = flag_l1_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1949" *) index_l1_20 : index_l1_21;
  assign index_l2_11[1:0] = flag_l1_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1950" *) index_l1_22 : index_l1_23;
  assign index_l2_12[1:0] = flag_l1_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1951" *) index_l1_24 : index_l1_25;
  assign index_l2_13[1:0] = flag_l1_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1952" *) index_l1_26 : index_l1_27;
  assign index_l2_14[1:0] = flag_l1_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1953" *) index_l1_28 : index_l1_29;
  assign index_l2_15[1:0] = flag_l1_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1954" *) index_l1_30 : index_l1_31;
  assign index_l2_16[1:0] = flag_l1_32 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1955" *) index_l1_32 : index_l1_33;
  assign index_l2_17[1:0] = flag_l1_34 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1956" *) index_l1_34 : index_l1_35;
  assign index_l2_18[1:0] = flag_l1_36 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1957" *) index_l1_36 : index_l1_37;
  assign index_l2_19[1:0] = flag_l1_38 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1958" *) index_l1_38 : index_l1_39;
  assign index_l2_20[1:0] = flag_l1_40 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1959" *) index_l1_40 : index_l1_41;
  assign index_l2_21[1:0] = flag_l1_42 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1960" *) index_l1_42 : index_l1_43;
  assign index_l2_22[1:0] = flag_l1_44 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1961" *) index_l1_44 : index_l1_45;
  assign index_l2_23[1:0] = flag_l1_46 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1962" *) index_l1_46 : index_l1_47;
  assign index_l2_24[1:0] = flag_l1_48 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1963" *) index_l1_48 : index_l1_49;
  assign index_l2_25[1:0] = flag_l1_50 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1964" *) index_l1_50 : index_l1_51;
  assign index_l2_26[1:0] = flag_l1_52 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1965" *) index_l1_52 : index_l1_53;
  assign index_l2_27[1:0] = flag_l1_54 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1966" *) index_l1_54 : index_l1_55;
  assign index_l2_28[1:0] = flag_l1_56 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1967" *) index_l1_56 : index_l1_57;
  assign index_l2_29[1:0] = flag_l1_58 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1968" *) index_l1_58 : index_l1_59;
  assign index_l2_30[1:0] = flag_l1_60 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1969" *) index_l1_60 : index_l1_61;
  assign index_l2_31[1:0] = flag_l1_62 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1970" *) index_l1_62 : index_l1_63;
  assign index_l3_0[2:0] = flag_l2_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1971" *) index_l2_0 : index_l2_1;
  assign index_l3_1[2:0] = flag_l2_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1972" *) index_l2_2 : index_l2_3;
  assign index_l3_2[2:0] = flag_l2_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1973" *) index_l2_4 : index_l2_5;
  assign index_l3_3[2:0] = flag_l2_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1974" *) index_l2_6 : index_l2_7;
  assign index_l3_4[2:0] = flag_l2_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1975" *) index_l2_8 : index_l2_9;
  assign index_l3_5[2:0] = flag_l2_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1976" *) index_l2_10 : index_l2_11;
  assign index_l3_6[2:0] = flag_l2_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1977" *) index_l2_12 : index_l2_13;
  assign index_l3_7[2:0] = flag_l2_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1978" *) index_l2_14 : index_l2_15;
  assign index_l3_8[2:0] = flag_l2_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1979" *) index_l2_16 : index_l2_17;
  assign index_l3_9[2:0] = flag_l2_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1980" *) index_l2_18 : index_l2_19;
  assign index_l3_10[2:0] = flag_l2_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1981" *) index_l2_20 : index_l2_21;
  assign index_l3_11[2:0] = flag_l2_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1982" *) index_l2_22 : index_l2_23;
  assign index_l3_12[2:0] = flag_l2_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1983" *) index_l2_24 : index_l2_25;
  assign index_l3_13[2:0] = flag_l2_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1984" *) index_l2_26 : index_l2_27;
  assign index_l3_14[2:0] = flag_l2_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1985" *) index_l2_28 : index_l2_29;
  assign index_l3_15[2:0] = flag_l2_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1986" *) index_l2_30 : index_l2_31;
  assign index_l4_0[3:0] = flag_l3_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1987" *) index_l3_0 : index_l3_1;
  assign index_l4_1[3:0] = flag_l3_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1988" *) index_l3_2 : index_l3_3;
  assign index_l4_2[3:0] = flag_l3_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1989" *) index_l3_4 : index_l3_5;
  assign index_l4_3[3:0] = flag_l3_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1990" *) index_l3_6 : index_l3_7;
  assign index_l4_4[3:0] = flag_l3_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1991" *) index_l3_8 : index_l3_9;
  assign index_l4_5[3:0] = flag_l3_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1992" *) index_l3_10 : index_l3_11;
  assign index_l4_6[3:0] = flag_l3_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1993" *) index_l3_12 : index_l3_13;
  assign index_l4_7[3:0] = flag_l3_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1994" *) index_l3_14 : index_l3_15;
  assign index_l5_0[4:0] = flag_l4_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1995" *) index_l4_0 : index_l4_1;
  assign index_l5_1[4:0] = flag_l4_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1996" *) index_l4_2 : index_l4_3;
  assign index_l5_2[4:0] = flag_l4_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1997" *) index_l4_4 : index_l4_5;
  assign index_l5_3[4:0] = flag_l4_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1998" *) index_l4_6 : index_l4_7;
  assign index_l6_0[5:0] = flag_l5_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:1999" *) index_l5_0 : index_l5_1;
  assign index_l6_1[5:0] = flag_l5_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2000" *) index_l5_2 : index_l5_3;
  assign adr_ram_wr_data[6:0] = flag_l6_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2001" *) index_l6_0 : index_l6_1;
  assign _2541_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2114" *) cq_rd_count0 : _0374_;
  assign _2542_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2115" *) _2531_ : cq_rd_count0;
  assign rd_count0_next = rd_pushing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2115" *) _2541_ : _2542_;
  assign _2543_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2117" *) cq_rd_count1 : _0375_;
  assign _2544_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2118" *) _2532_ : cq_rd_count1;
  assign rd_count1_next = rd_pushing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2118" *) _2543_ : _2544_;
  assign _2545_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2120" *) cq_rd_count2 : _0376_;
  assign _2546_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2121" *) _2533_ : cq_rd_count2;
  assign rd_count2_next = rd_pushing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2121" *) _2545_ : _2546_;
  assign _2547_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2123" *) cq_rd_count3 : _0377_;
  assign _2548_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2124" *) _2534_ : cq_rd_count3;
  assign rd_count3_next = rd_pushing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2124" *) _2547_ : _2548_;
  assign _2549_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2126" *) cq_rd_count4 : _0378_;
  assign _2550_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2127" *) _2535_ : cq_rd_count4;
  assign rd_count4_next = rd_pushing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2127" *) _2549_ : _2550_;
  assign _2551_ = rd_take5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2129" *) cq_rd_count5 : _0379_;
  assign _2552_ = rd_take5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2130" *) _2536_ : cq_rd_count5;
  assign rd_count5_next = rd_pushing5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2130" *) _2551_ : _2552_;
  assign _2553_ = rd_take6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2132" *) cq_rd_count6 : _0380_;
  assign _2554_ = rd_take6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2133" *) _2537_ : cq_rd_count6;
  assign rd_count6_next = rd_pushing6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2133" *) _2553_ : _2554_;
  assign _2555_ = rd_take7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2135" *) cq_rd_count7 : _0381_;
  assign _2556_ = rd_take7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2136" *) _2538_ : cq_rd_count7;
  assign rd_count7_next = rd_pushing7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2136" *) _2555_ : _2556_;
  assign _2557_ = rd_take8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2138" *) cq_rd_count8 : _0382_;
  assign _2558_ = rd_take8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2139" *) _2539_ : cq_rd_count8;
  assign rd_count8_next = rd_pushing8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2139" *) _2557_ : _2558_;
  assign _2559_ = rd_take9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2141" *) cq_rd_count9 : _0383_;
  assign _2560_ = rd_take9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2142" *) _2540_ : cq_rd_count9;
  assign rd_count9_next = rd_pushing9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2142" *) _2559_ : _2560_;
  assign _2561_ = _1224_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2491" *) adr_ram_rd_data : head0;
  assign _2562_ = _1225_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2492" *) adr_ram_rd_data : head1;
  assign _2563_ = _1226_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2493" *) adr_ram_rd_data : head2;
  assign _2564_ = _1227_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2494" *) adr_ram_rd_data : head3;
  assign _2565_ = _1228_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2495" *) adr_ram_rd_data : head4;
  assign _2566_ = _1229_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2496" *) adr_ram_rd_data : head5;
  assign _2567_ = _1230_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2497" *) adr_ram_rd_data : head6;
  assign _2568_ = _1231_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2498" *) adr_ram_rd_data : head7;
  assign _2569_ = _1232_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2499" *) adr_ram_rd_data : head8;
  assign _2570_ = _1233_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2500" *) adr_ram_rd_data : head9;
  assign cq_rd0_pd = rd_skid0_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2567" *) rd_skid0_0 : cq_wr_pd;
  assign _2571_ = rd_take_n_dly[0] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2570" *) cq_rd_pd_p : cq_wr_pd;
  assign _2572_ = rd_bypassing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2582" *) cq_wr_pd : cq_rd_pd_p;
  assign _0047_ = _1237_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2609" *) _2248_ : _2250_;
  assign _0049_ = _1237_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2610" *) _2251_ : _2252_;
  assign _0051_ = _1237_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2612" *) _1251_ : _2251_;
  assign cq_rd0_credits_next = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2621" *) cq_rd0_credits_w_take_next : cq_rd0_credits_wo_take_next;
  assign _2573_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2635" *) _2457_ : _2458_;
  assign cq_rd1_pd = rd_skid1_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2663" *) rd_skid1_0 : cq_wr_pd;
  assign _2574_ = rd_take_n_dly[1] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2666" *) cq_rd_pd_p : cq_wr_pd;
  assign _2575_ = rd_bypassing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2678" *) cq_wr_pd : cq_rd_pd_p;
  assign _0053_ = _1261_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2705" *) _2265_ : _2267_;
  assign _0055_ = _1261_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2706" *) _2268_ : _2269_;
  assign _0057_ = _1261_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2708" *) _1274_ : _2268_;
  assign cq_rd1_credits_next = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2717" *) cq_rd1_credits_w_take_next : cq_rd1_credits_wo_take_next;
  assign _2576_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2731" *) _2459_ : _2460_;
  assign cq_rd2_pd = rd_skid2_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2759" *) rd_skid2_0 : cq_wr_pd;
  assign _2577_ = rd_take_n_dly[2] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2762" *) cq_rd_pd_p : cq_wr_pd;
  assign _2578_ = rd_bypassing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2774" *) cq_wr_pd : cq_rd_pd_p;
  assign _0059_ = _1285_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2801" *) _2282_ : _2284_;
  assign _0061_ = _1285_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2802" *) _2285_ : _2286_;
  assign _0063_ = _1285_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2804" *) _1298_ : _2285_;
  assign cq_rd2_credits_next = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2813" *) cq_rd2_credits_w_take_next : cq_rd2_credits_wo_take_next;
  assign _2579_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2827" *) _2461_ : _2462_;
  assign cq_rd3_pd = rd_skid3_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2855" *) rd_skid3_0 : cq_wr_pd;
  assign _2580_ = rd_take_n_dly[3] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2858" *) cq_rd_pd_p : cq_wr_pd;
  assign _2581_ = rd_bypassing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2870" *) cq_wr_pd : cq_rd_pd_p;
  assign _0065_ = _1308_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2897" *) _2299_ : _2301_;
  assign _0067_ = _1308_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2898" *) _2302_ : _2303_;
  assign _0069_ = _1308_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2900" *) _1322_ : _2302_;
  assign cq_rd3_credits_next = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2909" *) cq_rd3_credits_w_take_next : cq_rd3_credits_wo_take_next;
  assign _2582_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2923" *) _2463_ : _2464_;
  assign cq_rd4_pd = rd_skid4_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2951" *) rd_skid4_0 : cq_wr_pd;
  assign _2583_ = rd_take_n_dly[4] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2954" *) cq_rd_pd_p : cq_wr_pd;
  assign _2584_ = rd_bypassing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2966" *) cq_wr_pd : cq_rd_pd_p;
  assign _0071_ = _1332_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2993" *) _2316_ : _2318_;
  assign _0073_ = _1332_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2994" *) _2319_ : _2320_;
  assign _0075_ = _1332_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2996" *) _1346_ : _2319_;
  assign cq_rd4_credits_next = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3005" *) cq_rd4_credits_w_take_next : cq_rd4_credits_wo_take_next;
  assign _2585_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3019" *) _2465_ : _2466_;
  assign cq_rd5_pd = rd_skid5_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3047" *) rd_skid5_0 : cq_wr_pd;
  assign _2586_ = rd_take_n_dly[5] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3050" *) cq_rd_pd_p : cq_wr_pd;
  assign _2587_ = rd_bypassing5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3062" *) cq_wr_pd : cq_rd_pd_p;
  assign _0077_ = _1356_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3089" *) _2333_ : _2335_;
  assign _0079_ = _1356_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3090" *) _2336_ : _2337_;
  assign _0081_ = _1356_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3092" *) _1370_ : _2336_;
  assign cq_rd5_credits_next = rd_take5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3101" *) cq_rd5_credits_w_take_next : cq_rd5_credits_wo_take_next;
  assign _2588_ = rd_take5 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3115" *) _2467_ : _2468_;
  assign cq_rd6_pd = rd_skid6_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3143" *) rd_skid6_0 : cq_wr_pd;
  assign _2589_ = rd_take_n_dly[6] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3146" *) cq_rd_pd_p : cq_wr_pd;
  assign _2590_ = rd_bypassing6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3158" *) cq_wr_pd : cq_rd_pd_p;
  assign _0083_ = _1380_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3185" *) _2350_ : _2352_;
  assign _0085_ = _1380_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3186" *) _2353_ : _2354_;
  assign _0087_ = _1380_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3188" *) _1393_ : _2353_;
  assign cq_rd6_credits_next = rd_take6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3197" *) cq_rd6_credits_w_take_next : cq_rd6_credits_wo_take_next;
  assign _2591_ = rd_take6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3211" *) _2469_ : _2470_;
  assign cq_rd7_pd = rd_skid7_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3239" *) rd_skid7_0 : cq_wr_pd;
  assign _2592_ = rd_take_n_dly[7] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3242" *) cq_rd_pd_p : cq_wr_pd;
  assign _2593_ = rd_bypassing7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3254" *) cq_wr_pd : cq_rd_pd_p;
  assign _0089_ = _1404_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3281" *) _2367_ : _2369_;
  assign _0091_ = _1404_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3282" *) _2370_ : _2371_;
  assign _0093_ = _1404_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3284" *) _1417_ : _2370_;
  assign cq_rd7_credits_next = rd_take7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3293" *) cq_rd7_credits_w_take_next : cq_rd7_credits_wo_take_next;
  assign _2594_ = rd_take7 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3307" *) _2471_ : _2472_;
  assign cq_rd8_pd = rd_skid8_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3335" *) rd_skid8_0 : cq_wr_pd;
  assign _2595_ = rd_take_n_dly[8] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3338" *) cq_rd_pd_p : cq_wr_pd;
  assign _2596_ = rd_bypassing8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3350" *) cq_wr_pd : cq_rd_pd_p;
  assign _0095_ = _1427_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3377" *) _2384_ : _2386_;
  assign _0097_ = _1427_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3378" *) _2387_ : _2388_;
  assign _0099_ = _1427_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3380" *) _1441_ : _2387_;
  assign cq_rd8_credits_next = rd_take8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3389" *) cq_rd8_credits_w_take_next : cq_rd8_credits_wo_take_next;
  assign _2597_ = rd_take8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3403" *) _2473_ : _2474_;
  assign cq_rd9_pd = rd_skid9_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3431" *) rd_skid9_0 : cq_wr_pd;
  assign _2598_ = rd_take_n_dly[9] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3434" *) cq_rd_pd_p : cq_wr_pd;
  assign _2599_ = rd_bypassing9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3446" *) cq_wr_pd : cq_rd_pd_p;
  assign _0101_ = _1451_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3473" *) _2401_ : _2403_;
  assign _0103_ = _1451_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3474" *) _2404_ : _2405_;
  assign _0105_ = _1451_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3476" *) _1465_ : _2404_;
  assign cq_rd9_credits_next = rd_take9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3485" *) cq_rd9_credits_w_take_next : cq_rd9_credits_wo_take_next;
  assign _2600_ = rd_take9 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:3499" *) _2475_ : _2476_;
  assign _2529_ = rd_pushing ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:162" *) rd_take_dly;
  assign _2528_ = rd_pushing0 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2156" *) rd_take0;
  assign _2527_ = rd_pushing1 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2165" *) rd_take1;
  assign _2526_ = rd_pushing2 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2174" *) rd_take2;
  assign _2525_ = rd_pushing3 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2183" *) rd_take3;
  assign _2524_ = rd_pushing4 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2192" *) rd_take4;
  assign _2523_ = rd_pushing5 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2201" *) rd_take5;
  assign _2522_ = rd_pushing6 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2210" *) rd_take6;
  assign _2521_ = rd_pushing7 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2219" *) rd_take7;
  assign _2520_ = rd_pushing8 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2228" *) rd_take8;
  assign _2519_ = rd_pushing9 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2237" *) rd_take9;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:2427" *)
  nv_ram_rwst_256x8 adr_ram (
    .clk(nvdla_core_clk),
    .di(adr_ram_wr_data),
    .dout(adr_ram_rd_data),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(adr_ram_rd_adr),
    .re(adr_ram_rd_enable),
    .wa(adr_ram_wr_adr),
    .we(adr_ram_wr_enable)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:108" *)
  NV_CLK_gate_power nvdla_core_clk_mgate (
    .clk(nvdla_core_clk),
    .clk_en(nvdla_core_clk_mgated_enable),
    .clk_gated(nvdla_core_clk_mgated),
    .reset_(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:105" *)
  NV_CLK_gate_power nvdla_core_clk_rd_mgate_skid (
    .clk(nvdla_core_clk),
    .clk_en(nvdla_core_clk_mgated_skid_enable),
    .clk_gated(nvdla_core_clk_mgated_skid),
    .reset_(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_MCIF_READ_cq.v:184" *)
  \$paramod\nv_ram_rws_256x7\FORCE_CONTENTION_ASSERTION_RESET_ACTIVE=1'1  ram (
    .clk(nvdla_core_clk),
    .di(cq_wr_pd),
    .dout(cq_rd_pd_p),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(adr_ram_rd_adr),
    .re(cq_rd_take),
    .wa(adr_ram_wr_data),
    .we(rd_pushing)
  );
  assign cq_rd_adr = adr_ram_rd_adr;
  assign cq_rd_adr_p = adr_ram_rd_adr;
  assign cq_wr_adr = adr_ram_wr_data;
  assign free_adr_index = adr_ram_wr_data;
  assign index_l7_0 = adr_ram_wr_data;
  assign rd_enable = cq_rd_take;
  assign rd_popping = rd_take_dly;
  assign rd_popping_adr = rd_adr_dly;
  assign rd_pushing_adr = adr_ram_wr_data;
  assign rd_pushing_thread_id = cq_wr_thread_id;
  assign rd_take_dly_cg = rd_take_dly;
  assign wr_adr_popping = rd_pushing;
  assign wr_count_next_is_256 = cq_wr_busy_next;
  assign wr_limit_muxed = 9'b000000000;
  assign wr_limit_reg = 9'b000000000;
  assign wr_popping = rd_take_dly;
  assign wr_pushing = rd_pushing;
  assign wr_pushing_thread_id = cq_wr_thread_id;
  assign wr_reserving_and_not_bypassing = rd_pushing;
endmodule
