module FP32_MUL_chn_b_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_mul.v:85" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_mul.v:86" *)
  output outsig;
  assign outsig = in_0;
endmodule
