module SDP_C_chn_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:329" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:330" *)
  output outsig;
  assign outsig = in_0;
endmodule
