module NV_NVDLA_CSC_WL_dec(nvdla_core_clk, nvdla_core_rstn, input_data, input_mask, input_mask_en, input_pipe_valid, input_sel, is_fp16, is_int8, output_data0, output_data1, output_data10, output_data100, output_data101, output_data102, output_data103, output_data104, output_data105, output_data106, output_data107, output_data108, output_data109, output_data11, output_data110, output_data111, output_data112, output_data113, output_data114, output_data115, output_data116, output_data117, output_data118, output_data119, output_data12, output_data120, output_data121, output_data122, output_data123, output_data124, output_data125, output_data126, output_data127, output_data13, output_data14, output_data15, output_data16, output_data17, output_data18, output_data19, output_data2, output_data20, output_data21, output_data22, output_data23, output_data24, output_data25, output_data26, output_data27, output_data28, output_data29, output_data3, output_data30, output_data31, output_data32, output_data33, output_data34, output_data35, output_data36, output_data37, output_data38, output_data39, output_data4, output_data40, output_data41, output_data42, output_data43, output_data44, output_data45, output_data46, output_data47, output_data48, output_data49, output_data5, output_data50, output_data51, output_data52, output_data53, output_data54, output_data55, output_data56, output_data57, output_data58, output_data59, output_data6, output_data60, output_data61, output_data62, output_data63, output_data64, output_data65, output_data66, output_data67, output_data68, output_data69, output_data7, output_data70, output_data71, output_data72, output_data73, output_data74, output_data75, output_data76, output_data77, output_data78, output_data79, output_data8, output_data80, output_data81, output_data82, output_data83, output_data84, output_data85, output_data86, output_data87, output_data88, output_data89, output_data9, output_data90, output_data91, output_data92, output_data93, output_data94, output_data95, output_data96, output_data97, output_data98, output_data99, output_mask, output_pvld, output_sel);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2575" *)
  wire [1023:0] _00000_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2585" *)
  wire [127:0] _00001_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21148" *)
  wire [127:0] _00002_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2595" *)
  wire [15:0] _00003_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13174" *)
  wire [15:0] _00004_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21158" *)
  wire [15:0] _00005_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13184" *)
  wire [7:0] _00006_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21168" *)
  wire [7:0] _00007_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13194" *)
  wire [7:0] _00008_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21178" *)
  wire [7:0] _00009_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13204" *)
  wire [7:0] _00010_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21188" *)
  wire [7:0] _00011_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13214" *)
  wire [7:0] _00012_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21198" *)
  wire [7:0] _00013_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13224" *)
  wire [7:0] _00014_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21208" *)
  wire [7:0] _00015_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13234" *)
  wire [7:0] _00016_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21218" *)
  wire [7:0] _00017_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13244" *)
  wire [7:0] _00018_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21228" *)
  wire [7:0] _00019_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13254" *)
  wire [7:0] _00020_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21238" *)
  wire [7:0] _00021_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13264" *)
  wire [7:0] _00022_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21248" *)
  wire [7:0] _00023_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13274" *)
  wire [7:0] _00024_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21258" *)
  wire [7:0] _00025_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13284" *)
  wire [7:0] _00026_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21268" *)
  wire [7:0] _00027_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13294" *)
  wire [7:0] _00028_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21278" *)
  wire [7:0] _00029_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13304" *)
  wire [7:0] _00030_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21288" *)
  wire [7:0] _00031_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13314" *)
  wire [7:0] _00032_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21298" *)
  wire [7:0] _00033_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13324" *)
  wire [7:0] _00034_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21308" *)
  wire [7:0] _00035_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13334" *)
  wire [7:0] _00036_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21318" *)
  wire [7:0] _00037_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13344" *)
  wire [7:0] _00038_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21328" *)
  wire [7:0] _00039_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13354" *)
  wire [7:0] _00040_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21338" *)
  wire [7:0] _00041_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13364" *)
  wire [7:0] _00042_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21348" *)
  wire [7:0] _00043_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13374" *)
  wire [7:0] _00044_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21358" *)
  wire [7:0] _00045_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13384" *)
  wire [7:0] _00046_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21368" *)
  wire [7:0] _00047_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13394" *)
  wire [7:0] _00048_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21378" *)
  wire [7:0] _00049_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13404" *)
  wire [7:0] _00050_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21388" *)
  wire [7:0] _00051_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13414" *)
  wire [7:0] _00052_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21398" *)
  wire [7:0] _00053_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13424" *)
  wire [7:0] _00054_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21408" *)
  wire [7:0] _00055_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13434" *)
  wire [7:0] _00056_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21418" *)
  wire [7:0] _00057_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13444" *)
  wire [7:0] _00058_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21428" *)
  wire [7:0] _00059_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13454" *)
  wire [7:0] _00060_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21438" *)
  wire [7:0] _00061_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13464" *)
  wire [7:0] _00062_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21448" *)
  wire [7:0] _00063_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13474" *)
  wire [7:0] _00064_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21458" *)
  wire [7:0] _00065_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13484" *)
  wire [7:0] _00066_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21468" *)
  wire [7:0] _00067_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13494" *)
  wire [7:0] _00068_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21478" *)
  wire [7:0] _00069_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13504" *)
  wire [7:0] _00070_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21488" *)
  wire [7:0] _00071_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13514" *)
  wire [7:0] _00072_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21498" *)
  wire [7:0] _00073_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13524" *)
  wire [7:0] _00074_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21508" *)
  wire [7:0] _00075_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13534" *)
  wire [7:0] _00076_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21518" *)
  wire [7:0] _00077_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13544" *)
  wire [7:0] _00078_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21528" *)
  wire [7:0] _00079_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13554" *)
  wire [7:0] _00080_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21538" *)
  wire [7:0] _00081_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13564" *)
  wire [7:0] _00082_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21548" *)
  wire [7:0] _00083_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13574" *)
  wire [7:0] _00084_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21558" *)
  wire [7:0] _00085_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13584" *)
  wire [7:0] _00086_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21568" *)
  wire [7:0] _00087_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13594" *)
  wire [7:0] _00088_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21578" *)
  wire [7:0] _00089_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13604" *)
  wire [7:0] _00090_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21588" *)
  wire [7:0] _00091_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13614" *)
  wire [7:0] _00092_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21598" *)
  wire [7:0] _00093_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13624" *)
  wire [7:0] _00094_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21608" *)
  wire [7:0] _00095_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13634" *)
  wire [7:0] _00096_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21618" *)
  wire [7:0] _00097_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13644" *)
  wire [7:0] _00098_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21628" *)
  wire [7:0] _00099_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13654" *)
  wire [7:0] _00100_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21638" *)
  wire [7:0] _00101_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13664" *)
  wire [7:0] _00102_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21648" *)
  wire [7:0] _00103_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13674" *)
  wire [7:0] _00104_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21658" *)
  wire [7:0] _00105_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13684" *)
  wire [7:0] _00106_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21668" *)
  wire [7:0] _00107_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13694" *)
  wire [7:0] _00108_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21678" *)
  wire [7:0] _00109_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13704" *)
  wire [7:0] _00110_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21688" *)
  wire [7:0] _00111_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13714" *)
  wire [7:0] _00112_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21698" *)
  wire [7:0] _00113_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13724" *)
  wire [7:0] _00114_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21708" *)
  wire [7:0] _00115_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13734" *)
  wire [7:0] _00116_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21718" *)
  wire [7:0] _00117_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13744" *)
  wire [7:0] _00118_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21728" *)
  wire [7:0] _00119_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13754" *)
  wire [7:0] _00120_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21738" *)
  wire [7:0] _00121_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13764" *)
  wire [7:0] _00122_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21748" *)
  wire [7:0] _00123_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13774" *)
  wire [7:0] _00124_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21758" *)
  wire [7:0] _00125_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13784" *)
  wire [7:0] _00126_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21768" *)
  wire [7:0] _00127_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13794" *)
  wire [7:0] _00128_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21778" *)
  wire [7:0] _00129_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13804" *)
  wire [7:0] _00130_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21788" *)
  wire [7:0] _00131_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13814" *)
  wire [7:0] _00132_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21798" *)
  wire [7:0] _00133_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13824" *)
  wire [7:0] _00134_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21808" *)
  wire [7:0] _00135_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13834" *)
  wire [7:0] _00136_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21818" *)
  wire [7:0] _00137_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13844" *)
  wire [7:0] _00138_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21828" *)
  wire [7:0] _00139_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13854" *)
  wire [7:0] _00140_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21838" *)
  wire [7:0] _00141_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13864" *)
  wire [7:0] _00142_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21848" *)
  wire [7:0] _00143_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13874" *)
  wire [7:0] _00144_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21858" *)
  wire [7:0] _00145_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13884" *)
  wire [7:0] _00146_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21868" *)
  wire [7:0] _00147_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13894" *)
  wire [7:0] _00148_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21878" *)
  wire [7:0] _00149_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13904" *)
  wire [7:0] _00150_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21888" *)
  wire [7:0] _00151_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13914" *)
  wire [7:0] _00152_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21898" *)
  wire [7:0] _00153_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13924" *)
  wire [7:0] _00154_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21908" *)
  wire [7:0] _00155_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13934" *)
  wire [7:0] _00156_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21918" *)
  wire [7:0] _00157_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13944" *)
  wire [7:0] _00158_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21928" *)
  wire [7:0] _00159_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13954" *)
  wire [7:0] _00160_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21938" *)
  wire [7:0] _00161_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13964" *)
  wire [7:0] _00162_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21948" *)
  wire [7:0] _00163_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13974" *)
  wire [7:0] _00164_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21958" *)
  wire [7:0] _00165_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13984" *)
  wire [7:0] _00166_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21968" *)
  wire [7:0] _00167_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13994" *)
  wire [7:0] _00168_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21978" *)
  wire [7:0] _00169_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14004" *)
  wire [7:0] _00170_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21988" *)
  wire [7:0] _00171_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14014" *)
  wire [7:0] _00172_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21998" *)
  wire [7:0] _00173_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14024" *)
  wire [7:0] _00174_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22008" *)
  wire [7:0] _00175_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14034" *)
  wire [7:0] _00176_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22018" *)
  wire [7:0] _00177_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14044" *)
  wire [7:0] _00178_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22028" *)
  wire [7:0] _00179_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14054" *)
  wire [7:0] _00180_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22038" *)
  wire [7:0] _00181_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14064" *)
  wire [7:0] _00182_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22048" *)
  wire [7:0] _00183_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14074" *)
  wire [7:0] _00184_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22058" *)
  wire [7:0] _00185_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14084" *)
  wire [7:0] _00186_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22068" *)
  wire [7:0] _00187_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14094" *)
  wire [7:0] _00188_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22078" *)
  wire [7:0] _00189_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14104" *)
  wire [7:0] _00190_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22088" *)
  wire [7:0] _00191_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14114" *)
  wire [7:0] _00192_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22098" *)
  wire [7:0] _00193_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14124" *)
  wire [7:0] _00194_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22108" *)
  wire [7:0] _00195_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14134" *)
  wire [7:0] _00196_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22118" *)
  wire [7:0] _00197_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14144" *)
  wire [7:0] _00198_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22128" *)
  wire [7:0] _00199_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14154" *)
  wire [7:0] _00200_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22138" *)
  wire [7:0] _00201_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14164" *)
  wire [7:0] _00202_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22148" *)
  wire [7:0] _00203_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14174" *)
  wire [7:0] _00204_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22158" *)
  wire [7:0] _00205_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14184" *)
  wire [7:0] _00206_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22168" *)
  wire [7:0] _00207_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14194" *)
  wire [7:0] _00208_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22178" *)
  wire [7:0] _00209_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14204" *)
  wire [7:0] _00210_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22188" *)
  wire [7:0] _00211_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14214" *)
  wire [7:0] _00212_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22198" *)
  wire [7:0] _00213_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14224" *)
  wire [7:0] _00214_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22208" *)
  wire [7:0] _00215_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14234" *)
  wire [7:0] _00216_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22218" *)
  wire [7:0] _00217_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14244" *)
  wire [7:0] _00218_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22228" *)
  wire [7:0] _00219_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14254" *)
  wire [7:0] _00220_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22238" *)
  wire [7:0] _00221_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14264" *)
  wire [7:0] _00222_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22248" *)
  wire [7:0] _00223_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14274" *)
  wire [7:0] _00224_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22258" *)
  wire [7:0] _00225_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14284" *)
  wire [7:0] _00226_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22268" *)
  wire [7:0] _00227_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14294" *)
  wire [7:0] _00228_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22278" *)
  wire [7:0] _00229_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14304" *)
  wire [7:0] _00230_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22288" *)
  wire [7:0] _00231_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14314" *)
  wire [7:0] _00232_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22298" *)
  wire [7:0] _00233_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14324" *)
  wire [7:0] _00234_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22308" *)
  wire [7:0] _00235_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14334" *)
  wire [7:0] _00236_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22318" *)
  wire [7:0] _00237_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14344" *)
  wire [7:0] _00238_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22328" *)
  wire [7:0] _00239_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14354" *)
  wire [7:0] _00240_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22338" *)
  wire [7:0] _00241_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14364" *)
  wire [7:0] _00242_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22348" *)
  wire [7:0] _00243_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14374" *)
  wire [7:0] _00244_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22358" *)
  wire [7:0] _00245_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14384" *)
  wire [7:0] _00246_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22368" *)
  wire [7:0] _00247_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14394" *)
  wire [7:0] _00248_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22378" *)
  wire [7:0] _00249_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14404" *)
  wire [7:0] _00250_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22388" *)
  wire [7:0] _00251_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14414" *)
  wire [7:0] _00252_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22398" *)
  wire [7:0] _00253_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14424" *)
  wire [7:0] _00254_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22408" *)
  wire [7:0] _00255_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14434" *)
  wire [7:0] _00256_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22418" *)
  wire [7:0] _00257_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14444" *)
  wire [7:0] _00258_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22428" *)
  wire [7:0] _00259_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14454" *)
  wire [7:0] _00260_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22438" *)
  wire [7:0] _00261_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2605" *)
  wire _00262_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2615" *)
  wire [1:0] _00263_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2625" *)
  wire [1:0] _00264_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2635" *)
  wire [2:0] _00265_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2645" *)
  wire [2:0] _00266_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2655" *)
  wire [2:0] _00267_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2665" *)
  wire [2:0] _00268_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2675" *)
  wire [3:0] _00269_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2685" *)
  wire [3:0] _00270_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2695" *)
  wire [3:0] _00271_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2705" *)
  wire [3:0] _00272_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2715" *)
  wire [3:0] _00273_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2725" *)
  wire [3:0] _00274_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2735" *)
  wire [3:0] _00275_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2745" *)
  wire [3:0] _00276_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2755" *)
  wire [4:0] _00277_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2765" *)
  wire [4:0] _00278_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2775" *)
  wire [4:0] _00279_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2785" *)
  wire [4:0] _00280_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2795" *)
  wire [4:0] _00281_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2805" *)
  wire [4:0] _00282_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2815" *)
  wire [4:0] _00283_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2825" *)
  wire [4:0] _00284_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2835" *)
  wire [4:0] _00285_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2845" *)
  wire [4:0] _00286_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2855" *)
  wire [4:0] _00287_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2865" *)
  wire [4:0] _00288_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2875" *)
  wire [4:0] _00289_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2885" *)
  wire [4:0] _00290_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2895" *)
  wire [4:0] _00291_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2905" *)
  wire [4:0] _00292_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2915" *)
  wire [5:0] _00293_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2925" *)
  wire [5:0] _00294_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2935" *)
  wire [5:0] _00295_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2945" *)
  wire [5:0] _00296_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2955" *)
  wire [5:0] _00297_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2965" *)
  wire [5:0] _00298_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2975" *)
  wire [5:0] _00299_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2985" *)
  wire [5:0] _00300_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2995" *)
  wire [5:0] _00301_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3005" *)
  wire [5:0] _00302_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3015" *)
  wire [5:0] _00303_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3025" *)
  wire [5:0] _00304_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3035" *)
  wire [5:0] _00305_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3045" *)
  wire [5:0] _00306_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3055" *)
  wire [5:0] _00307_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3065" *)
  wire [5:0] _00308_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3075" *)
  wire [5:0] _00309_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3085" *)
  wire [5:0] _00310_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3095" *)
  wire [5:0] _00311_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3105" *)
  wire [5:0] _00312_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3115" *)
  wire [5:0] _00313_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3125" *)
  wire [5:0] _00314_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3135" *)
  wire [5:0] _00315_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3145" *)
  wire [5:0] _00316_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3155" *)
  wire [5:0] _00317_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3165" *)
  wire [5:0] _00318_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3175" *)
  wire [5:0] _00319_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3185" *)
  wire [5:0] _00320_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3195" *)
  wire [5:0] _00321_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3205" *)
  wire [5:0] _00322_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3215" *)
  wire [5:0] _00323_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3225" *)
  wire [5:0] _00324_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3235" *)
  wire [6:0] _00325_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3245" *)
  wire [6:0] _00326_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3255" *)
  wire [6:0] _00327_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3265" *)
  wire [6:0] _00328_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3275" *)
  wire [6:0] _00329_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3285" *)
  wire [6:0] _00330_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3295" *)
  wire [6:0] _00331_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3305" *)
  wire [6:0] _00332_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3315" *)
  wire [6:0] _00333_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3325" *)
  wire [6:0] _00334_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3335" *)
  wire [6:0] _00335_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3345" *)
  wire [6:0] _00336_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3355" *)
  wire [6:0] _00337_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3365" *)
  wire [6:0] _00338_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3375" *)
  wire [6:0] _00339_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3385" *)
  wire [6:0] _00340_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3395" *)
  wire [6:0] _00341_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3405" *)
  wire [6:0] _00342_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3415" *)
  wire [6:0] _00343_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3425" *)
  wire [6:0] _00344_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3435" *)
  wire [6:0] _00345_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3445" *)
  wire [6:0] _00346_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3455" *)
  wire [6:0] _00347_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3465" *)
  wire [6:0] _00348_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3475" *)
  wire [6:0] _00349_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3485" *)
  wire [6:0] _00350_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3495" *)
  wire [6:0] _00351_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3505" *)
  wire [6:0] _00352_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3515" *)
  wire [6:0] _00353_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3525" *)
  wire [6:0] _00354_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3535" *)
  wire [6:0] _00355_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3545" *)
  wire [6:0] _00356_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3555" *)
  wire [6:0] _00357_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3565" *)
  wire [6:0] _00358_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3575" *)
  wire [6:0] _00359_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3585" *)
  wire [6:0] _00360_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3595" *)
  wire [6:0] _00361_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3605" *)
  wire [6:0] _00362_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3615" *)
  wire [6:0] _00363_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3625" *)
  wire [6:0] _00364_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3635" *)
  wire [6:0] _00365_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3645" *)
  wire [6:0] _00366_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3655" *)
  wire [6:0] _00367_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3665" *)
  wire [6:0] _00368_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3675" *)
  wire [6:0] _00369_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3685" *)
  wire [6:0] _00370_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3695" *)
  wire [6:0] _00371_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3705" *)
  wire [6:0] _00372_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3715" *)
  wire [6:0] _00373_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3725" *)
  wire [6:0] _00374_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3735" *)
  wire [6:0] _00375_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3745" *)
  wire [6:0] _00376_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3755" *)
  wire [6:0] _00377_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3765" *)
  wire [6:0] _00378_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3775" *)
  wire [6:0] _00379_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3785" *)
  wire [6:0] _00380_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3795" *)
  wire [6:0] _00381_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3805" *)
  wire [6:0] _00382_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3815" *)
  wire [6:0] _00383_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3825" *)
  wire [6:0] _00384_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3835" *)
  wire [6:0] _00385_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3845" *)
  wire [6:0] _00386_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3855" *)
  wire [6:0] _00387_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3865" *)
  wire [6:0] _00388_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3875" *)
  wire [7:0] _00389_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *)
  wire [2:0] _00390_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *)
  wire [3:0] _00391_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *)
  wire [3:0] _00392_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *)
  wire [3:0] _00393_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *)
  wire [3:0] _00394_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *)
  wire [4:0] _00395_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *)
  wire [4:0] _00396_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *)
  wire [4:0] _00397_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00398_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00399_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00400_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00401_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00402_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00403_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00404_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *)
  wire [4:0] _00405_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1170" *)
  wire [5:0] _00406_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1170" *)
  wire [5:0] _00407_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00408_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00409_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00410_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00411_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00412_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00413_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00414_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *)
  wire [5:0] _00415_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00416_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00417_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00418_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00419_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00420_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00421_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00422_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *)
  wire [5:0] _00423_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00424_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00425_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00426_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00427_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00428_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00429_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00430_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *)
  wire [5:0] _00431_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1502" *)
  wire [6:0] _00432_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00433_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00434_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00435_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00436_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00437_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00438_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00439_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *)
  wire [6:0] _00440_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00441_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00442_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00443_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00444_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00445_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00446_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00447_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *)
  wire [6:0] _00448_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00449_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00450_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00451_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00452_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00453_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00454_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00455_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *)
  wire [6:0] _00456_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00457_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00458_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00459_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00460_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00461_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00462_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00463_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *)
  wire [6:0] _00464_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00465_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00466_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00467_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00468_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00469_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00470_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00471_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *)
  wire [6:0] _00472_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00473_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00474_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00475_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00476_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00477_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00478_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00479_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *)
  wire [6:0] _00480_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00481_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00482_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00483_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00484_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00485_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00486_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00487_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *)
  wire [6:0] _00488_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00489_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00490_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00491_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00492_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00493_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00494_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00495_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *)
  wire [7:0] _00496_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00497_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00498_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00499_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00500_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00501_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00502_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00503_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *)
  wire [7:0] _00504_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00505_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00506_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00507_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00508_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00509_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00510_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00511_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *)
  wire [7:0] _00512_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00513_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00514_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00515_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00516_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00517_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00518_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00519_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *)
  wire [7:0] _00520_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00521_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00522_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00523_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00524_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00525_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00526_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00527_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *)
  wire [7:0] _00528_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00529_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00530_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00531_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00532_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00533_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00534_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00535_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *)
  wire [7:0] _00536_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00537_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00538_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00539_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00540_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00541_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00542_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00543_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *)
  wire [7:0] _00544_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00545_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00546_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00547_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00548_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00549_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00550_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00551_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *)
  wire [7:0] _00552_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00553_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00554_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00555_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00556_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00557_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00558_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00559_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *)
  wire [7:0] _00560_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00561_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00562_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00563_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00564_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00565_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00566_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00567_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *)
  wire [7:0] _00568_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00569_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00570_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00571_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00572_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00573_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00574_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00575_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *)
  wire [7:0] _00576_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00577_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00578_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00579_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00580_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00581_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00582_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00583_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *)
  wire [7:0] _00584_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00585_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00586_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00587_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00588_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00589_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00590_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00591_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *)
  wire [7:0] _00592_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00593_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00594_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00595_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00596_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00597_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00598_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00599_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *)
  wire [7:0] _00600_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00601_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00602_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00603_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00604_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00605_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00606_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00607_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *)
  wire [7:0] _00608_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13186" *)
  wire [7:0] _00609_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13196" *)
  wire [7:0] _00610_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13206" *)
  wire [7:0] _00611_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13216" *)
  wire [7:0] _00612_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13226" *)
  wire [7:0] _00613_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13236" *)
  wire [7:0] _00614_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13246" *)
  wire [7:0] _00615_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13256" *)
  wire [7:0] _00616_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13266" *)
  wire [7:0] _00617_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13276" *)
  wire [7:0] _00618_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13286" *)
  wire [7:0] _00619_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13296" *)
  wire [7:0] _00620_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13306" *)
  wire [7:0] _00621_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13316" *)
  wire [7:0] _00622_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13326" *)
  wire [7:0] _00623_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13336" *)
  wire [7:0] _00624_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13346" *)
  wire [7:0] _00625_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13356" *)
  wire [7:0] _00626_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13366" *)
  wire [7:0] _00627_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13376" *)
  wire [7:0] _00628_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13386" *)
  wire [7:0] _00629_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13396" *)
  wire [7:0] _00630_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13406" *)
  wire [7:0] _00631_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13416" *)
  wire [7:0] _00632_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13426" *)
  wire [7:0] _00633_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13436" *)
  wire [7:0] _00634_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13446" *)
  wire [7:0] _00635_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13456" *)
  wire [7:0] _00636_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13466" *)
  wire [7:0] _00637_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13476" *)
  wire [7:0] _00638_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13486" *)
  wire [7:0] _00639_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13496" *)
  wire [7:0] _00640_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13506" *)
  wire [7:0] _00641_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13516" *)
  wire [7:0] _00642_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13526" *)
  wire [7:0] _00643_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13536" *)
  wire [7:0] _00644_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13546" *)
  wire [7:0] _00645_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13556" *)
  wire [7:0] _00646_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13566" *)
  wire [7:0] _00647_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13576" *)
  wire [7:0] _00648_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13586" *)
  wire [7:0] _00649_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13596" *)
  wire [7:0] _00650_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13606" *)
  wire [7:0] _00651_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13616" *)
  wire [7:0] _00652_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13626" *)
  wire [7:0] _00653_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13636" *)
  wire [7:0] _00654_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13646" *)
  wire [7:0] _00655_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13656" *)
  wire [7:0] _00656_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13666" *)
  wire [7:0] _00657_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13676" *)
  wire [7:0] _00658_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13686" *)
  wire [7:0] _00659_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13696" *)
  wire [7:0] _00660_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13706" *)
  wire [7:0] _00661_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13716" *)
  wire [7:0] _00662_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13726" *)
  wire [7:0] _00663_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13736" *)
  wire [7:0] _00664_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13746" *)
  wire [7:0] _00665_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13756" *)
  wire [7:0] _00666_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13766" *)
  wire [7:0] _00667_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13776" *)
  wire [7:0] _00668_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13786" *)
  wire [7:0] _00669_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13796" *)
  wire [7:0] _00670_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13806" *)
  wire [7:0] _00671_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13816" *)
  wire [7:0] _00672_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13826" *)
  wire [7:0] _00673_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13836" *)
  wire [7:0] _00674_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13846" *)
  wire [7:0] _00675_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13856" *)
  wire [7:0] _00676_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13866" *)
  wire [7:0] _00677_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13876" *)
  wire [7:0] _00678_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13886" *)
  wire [7:0] _00679_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13896" *)
  wire [7:0] _00680_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13906" *)
  wire [7:0] _00681_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13916" *)
  wire [7:0] _00682_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13926" *)
  wire [7:0] _00683_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13936" *)
  wire [7:0] _00684_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13946" *)
  wire [7:0] _00685_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13956" *)
  wire [7:0] _00686_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13966" *)
  wire [7:0] _00687_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13976" *)
  wire [7:0] _00688_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13986" *)
  wire [7:0] _00689_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13996" *)
  wire [7:0] _00690_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14006" *)
  wire [7:0] _00691_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14016" *)
  wire [7:0] _00692_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14026" *)
  wire [7:0] _00693_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14036" *)
  wire [7:0] _00694_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14046" *)
  wire [7:0] _00695_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14056" *)
  wire [7:0] _00696_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14066" *)
  wire [7:0] _00697_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14076" *)
  wire [7:0] _00698_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14086" *)
  wire [7:0] _00699_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14096" *)
  wire [7:0] _00700_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14106" *)
  wire [7:0] _00701_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14116" *)
  wire [7:0] _00702_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14126" *)
  wire [7:0] _00703_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14136" *)
  wire [7:0] _00704_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14146" *)
  wire [7:0] _00705_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14156" *)
  wire [7:0] _00706_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14166" *)
  wire [7:0] _00707_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14176" *)
  wire [7:0] _00708_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14186" *)
  wire [7:0] _00709_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14196" *)
  wire [7:0] _00710_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14206" *)
  wire [7:0] _00711_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14216" *)
  wire [7:0] _00712_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14226" *)
  wire [7:0] _00713_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14236" *)
  wire [7:0] _00714_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14246" *)
  wire [7:0] _00715_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14256" *)
  wire [7:0] _00716_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14266" *)
  wire [7:0] _00717_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14276" *)
  wire [7:0] _00718_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14286" *)
  wire [7:0] _00719_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14296" *)
  wire [7:0] _00720_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14306" *)
  wire [7:0] _00721_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14316" *)
  wire [7:0] _00722_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14326" *)
  wire [7:0] _00723_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14336" *)
  wire [7:0] _00724_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14346" *)
  wire [7:0] _00725_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14356" *)
  wire [7:0] _00726_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14366" *)
  wire [7:0] _00727_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14376" *)
  wire [7:0] _00728_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14386" *)
  wire [7:0] _00729_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14396" *)
  wire [7:0] _00730_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14406" *)
  wire [7:0] _00731_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14416" *)
  wire [7:0] _00732_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14426" *)
  wire [7:0] _00733_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14436" *)
  wire [7:0] _00734_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14446" *)
  wire [7:0] _00735_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14456" *)
  wire [7:0] _00736_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2606" *)
  wire _00737_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2766" *)
  wire _00738_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2926" *)
  wire _00739_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3086" *)
  wire _00740_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3246" *)
  wire _00741_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3406" *)
  wire _00742_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3566" *)
  wire _00743_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3726" *)
  wire _00744_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:944" *)
  wire [7:0] _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21139" *)
  wire [127:0] _09001_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:292" *)
  reg [1023:0] data_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:153" *)
  input [1023:0] input_data;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:154" *)
  input [127:0] input_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:155" *)
  input [9:0] input_mask_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:291" *)
  wire [127:0] input_mask_gated;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:156" *)
  input input_pipe_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:157" *)
  input [15:0] input_sel;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:158" *)
  input is_fp16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:159" *)
  input is_int8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:293" *)
  reg [127:0] mask_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:294" *)
  wire [127:0] mask_d2_fp16_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:295" *)
  wire [127:0] mask_d2_int16_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:296" *)
  wire [127:0] mask_d2_int8_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:297" *)
  wire [127:0] mask_d2_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:298" *)
  reg [127:0] mask_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:151" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:152" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:160" *)
  output [7:0] output_data0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:161" *)
  output [7:0] output_data1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:162" *)
  output [7:0] output_data10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:163" *)
  output [7:0] output_data100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:164" *)
  output [7:0] output_data101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:165" *)
  output [7:0] output_data102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:166" *)
  output [7:0] output_data103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:167" *)
  output [7:0] output_data104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:168" *)
  output [7:0] output_data105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:169" *)
  output [7:0] output_data106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:170" *)
  output [7:0] output_data107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:171" *)
  output [7:0] output_data108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:172" *)
  output [7:0] output_data109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:173" *)
  output [7:0] output_data11;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:174" *)
  output [7:0] output_data110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:175" *)
  output [7:0] output_data111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:176" *)
  output [7:0] output_data112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:177" *)
  output [7:0] output_data113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:178" *)
  output [7:0] output_data114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:179" *)
  output [7:0] output_data115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:180" *)
  output [7:0] output_data116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:181" *)
  output [7:0] output_data117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:182" *)
  output [7:0] output_data118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:183" *)
  output [7:0] output_data119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:184" *)
  output [7:0] output_data12;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:185" *)
  output [7:0] output_data120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:186" *)
  output [7:0] output_data121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:187" *)
  output [7:0] output_data122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:188" *)
  output [7:0] output_data123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:189" *)
  output [7:0] output_data124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:190" *)
  output [7:0] output_data125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:191" *)
  output [7:0] output_data126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:192" *)
  output [7:0] output_data127;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:193" *)
  output [7:0] output_data13;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:194" *)
  output [7:0] output_data14;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:195" *)
  output [7:0] output_data15;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:196" *)
  output [7:0] output_data16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:197" *)
  output [7:0] output_data17;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:198" *)
  output [7:0] output_data18;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:199" *)
  output [7:0] output_data19;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:200" *)
  output [7:0] output_data2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:201" *)
  output [7:0] output_data20;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:202" *)
  output [7:0] output_data21;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:203" *)
  output [7:0] output_data22;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:204" *)
  output [7:0] output_data23;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:205" *)
  output [7:0] output_data24;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:206" *)
  output [7:0] output_data25;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:207" *)
  output [7:0] output_data26;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:208" *)
  output [7:0] output_data27;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:209" *)
  output [7:0] output_data28;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:210" *)
  output [7:0] output_data29;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:211" *)
  output [7:0] output_data3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:212" *)
  output [7:0] output_data30;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:213" *)
  output [7:0] output_data31;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:214" *)
  output [7:0] output_data32;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:215" *)
  output [7:0] output_data33;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:216" *)
  output [7:0] output_data34;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:217" *)
  output [7:0] output_data35;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:218" *)
  output [7:0] output_data36;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:219" *)
  output [7:0] output_data37;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:220" *)
  output [7:0] output_data38;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:221" *)
  output [7:0] output_data39;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:222" *)
  output [7:0] output_data4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:223" *)
  output [7:0] output_data40;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:224" *)
  output [7:0] output_data41;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:225" *)
  output [7:0] output_data42;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:226" *)
  output [7:0] output_data43;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:227" *)
  output [7:0] output_data44;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:228" *)
  output [7:0] output_data45;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:229" *)
  output [7:0] output_data46;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:230" *)
  output [7:0] output_data47;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:231" *)
  output [7:0] output_data48;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:232" *)
  output [7:0] output_data49;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:233" *)
  output [7:0] output_data5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:234" *)
  output [7:0] output_data50;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:235" *)
  output [7:0] output_data51;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:236" *)
  output [7:0] output_data52;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:237" *)
  output [7:0] output_data53;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:238" *)
  output [7:0] output_data54;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:239" *)
  output [7:0] output_data55;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:240" *)
  output [7:0] output_data56;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:241" *)
  output [7:0] output_data57;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:242" *)
  output [7:0] output_data58;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:243" *)
  output [7:0] output_data59;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:244" *)
  output [7:0] output_data6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:245" *)
  output [7:0] output_data60;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:246" *)
  output [7:0] output_data61;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:247" *)
  output [7:0] output_data62;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:248" *)
  output [7:0] output_data63;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:249" *)
  output [7:0] output_data64;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:250" *)
  output [7:0] output_data65;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:251" *)
  output [7:0] output_data66;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:252" *)
  output [7:0] output_data67;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:253" *)
  output [7:0] output_data68;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:254" *)
  output [7:0] output_data69;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:255" *)
  output [7:0] output_data7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:256" *)
  output [7:0] output_data70;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:257" *)
  output [7:0] output_data71;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:258" *)
  output [7:0] output_data72;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:259" *)
  output [7:0] output_data73;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:260" *)
  output [7:0] output_data74;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:261" *)
  output [7:0] output_data75;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:262" *)
  output [7:0] output_data76;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:263" *)
  output [7:0] output_data77;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:264" *)
  output [7:0] output_data78;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:265" *)
  output [7:0] output_data79;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:266" *)
  output [7:0] output_data8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:267" *)
  output [7:0] output_data80;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:268" *)
  output [7:0] output_data81;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:269" *)
  output [7:0] output_data82;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:270" *)
  output [7:0] output_data83;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:271" *)
  output [7:0] output_data84;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:272" *)
  output [7:0] output_data85;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:273" *)
  output [7:0] output_data86;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:274" *)
  output [7:0] output_data87;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:275" *)
  output [7:0] output_data88;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:276" *)
  output [7:0] output_data89;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:277" *)
  output [7:0] output_data9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:278" *)
  output [7:0] output_data90;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:279" *)
  output [7:0] output_data91;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:280" *)
  output [7:0] output_data92;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:281" *)
  output [7:0] output_data93;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:282" *)
  output [7:0] output_data94;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:283" *)
  output [7:0] output_data95;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:284" *)
  output [7:0] output_data96;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:285" *)
  output [7:0] output_data97;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:286" *)
  output [7:0] output_data98;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:287" *)
  output [7:0] output_data99;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:288" *)
  output [127:0] output_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:289" *)
  output output_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:290" *)
  output [15:0] output_sel;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:299" *)
  reg [15:0] sel_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:300" *)
  reg [15:0] sel_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:301" *)
  reg [15:0] sel_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:302" *)
  reg valid_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:303" *)
  reg valid_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:304" *)
  reg valid_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:305" *)
  wire [7:0] vec_data_000;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:306" *)
  reg [7:0] vec_data_000_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:307" *)
  reg [7:0] vec_data_000_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:308" *)
  wire [7:0] vec_data_001;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:309" *)
  reg [7:0] vec_data_001_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:310" *)
  reg [7:0] vec_data_001_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:311" *)
  wire [7:0] vec_data_002;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:312" *)
  reg [7:0] vec_data_002_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:313" *)
  reg [7:0] vec_data_002_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:314" *)
  wire [7:0] vec_data_003;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:315" *)
  reg [7:0] vec_data_003_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:316" *)
  reg [7:0] vec_data_003_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:317" *)
  wire [7:0] vec_data_004;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:318" *)
  reg [7:0] vec_data_004_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:319" *)
  reg [7:0] vec_data_004_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:320" *)
  wire [7:0] vec_data_005;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:321" *)
  reg [7:0] vec_data_005_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:322" *)
  reg [7:0] vec_data_005_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:323" *)
  wire [7:0] vec_data_006;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:324" *)
  reg [7:0] vec_data_006_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:325" *)
  reg [7:0] vec_data_006_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:326" *)
  wire [7:0] vec_data_007;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:327" *)
  reg [7:0] vec_data_007_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:328" *)
  reg [7:0] vec_data_007_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:329" *)
  wire [7:0] vec_data_008;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:330" *)
  reg [7:0] vec_data_008_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:331" *)
  reg [7:0] vec_data_008_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:332" *)
  wire [7:0] vec_data_009;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:333" *)
  reg [7:0] vec_data_009_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:334" *)
  reg [7:0] vec_data_009_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:335" *)
  wire [7:0] vec_data_010;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:336" *)
  reg [7:0] vec_data_010_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:337" *)
  reg [7:0] vec_data_010_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:338" *)
  wire [7:0] vec_data_011;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:339" *)
  reg [7:0] vec_data_011_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:340" *)
  reg [7:0] vec_data_011_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:341" *)
  wire [7:0] vec_data_012;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:342" *)
  reg [7:0] vec_data_012_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:343" *)
  reg [7:0] vec_data_012_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:344" *)
  wire [7:0] vec_data_013;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:345" *)
  reg [7:0] vec_data_013_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:346" *)
  reg [7:0] vec_data_013_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:347" *)
  wire [7:0] vec_data_014;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:348" *)
  reg [7:0] vec_data_014_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:349" *)
  reg [7:0] vec_data_014_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:350" *)
  wire [7:0] vec_data_015;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:351" *)
  reg [7:0] vec_data_015_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:352" *)
  reg [7:0] vec_data_015_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:353" *)
  wire [7:0] vec_data_016;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:354" *)
  reg [7:0] vec_data_016_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:355" *)
  reg [7:0] vec_data_016_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:356" *)
  wire [7:0] vec_data_017;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:357" *)
  reg [7:0] vec_data_017_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:358" *)
  reg [7:0] vec_data_017_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:359" *)
  wire [7:0] vec_data_018;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:360" *)
  reg [7:0] vec_data_018_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:361" *)
  reg [7:0] vec_data_018_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:362" *)
  wire [7:0] vec_data_019;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:363" *)
  reg [7:0] vec_data_019_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:364" *)
  reg [7:0] vec_data_019_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:365" *)
  wire [7:0] vec_data_020;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:366" *)
  reg [7:0] vec_data_020_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:367" *)
  reg [7:0] vec_data_020_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:368" *)
  wire [7:0] vec_data_021;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:369" *)
  reg [7:0] vec_data_021_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:370" *)
  reg [7:0] vec_data_021_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:371" *)
  wire [7:0] vec_data_022;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:372" *)
  reg [7:0] vec_data_022_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:373" *)
  reg [7:0] vec_data_022_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:374" *)
  wire [7:0] vec_data_023;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:375" *)
  reg [7:0] vec_data_023_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:376" *)
  reg [7:0] vec_data_023_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:377" *)
  wire [7:0] vec_data_024;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:378" *)
  reg [7:0] vec_data_024_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:379" *)
  reg [7:0] vec_data_024_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:380" *)
  wire [7:0] vec_data_025;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:381" *)
  reg [7:0] vec_data_025_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:382" *)
  reg [7:0] vec_data_025_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:383" *)
  wire [7:0] vec_data_026;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:384" *)
  reg [7:0] vec_data_026_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:385" *)
  reg [7:0] vec_data_026_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:386" *)
  wire [7:0] vec_data_027;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:387" *)
  reg [7:0] vec_data_027_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:388" *)
  reg [7:0] vec_data_027_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:389" *)
  wire [7:0] vec_data_028;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:390" *)
  reg [7:0] vec_data_028_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:391" *)
  reg [7:0] vec_data_028_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:392" *)
  wire [7:0] vec_data_029;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:393" *)
  reg [7:0] vec_data_029_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:394" *)
  reg [7:0] vec_data_029_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:395" *)
  wire [7:0] vec_data_030;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:396" *)
  reg [7:0] vec_data_030_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:397" *)
  reg [7:0] vec_data_030_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:398" *)
  wire [7:0] vec_data_031;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:399" *)
  reg [7:0] vec_data_031_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:400" *)
  reg [7:0] vec_data_031_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:401" *)
  wire [7:0] vec_data_032;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:402" *)
  reg [7:0] vec_data_032_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:403" *)
  reg [7:0] vec_data_032_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:404" *)
  wire [7:0] vec_data_033;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:405" *)
  reg [7:0] vec_data_033_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:406" *)
  reg [7:0] vec_data_033_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:407" *)
  wire [7:0] vec_data_034;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:408" *)
  reg [7:0] vec_data_034_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:409" *)
  reg [7:0] vec_data_034_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:410" *)
  wire [7:0] vec_data_035;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:411" *)
  reg [7:0] vec_data_035_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:412" *)
  reg [7:0] vec_data_035_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:413" *)
  wire [7:0] vec_data_036;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:414" *)
  reg [7:0] vec_data_036_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:415" *)
  reg [7:0] vec_data_036_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:416" *)
  wire [7:0] vec_data_037;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:417" *)
  reg [7:0] vec_data_037_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:418" *)
  reg [7:0] vec_data_037_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:419" *)
  wire [7:0] vec_data_038;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:420" *)
  reg [7:0] vec_data_038_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:421" *)
  reg [7:0] vec_data_038_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:422" *)
  wire [7:0] vec_data_039;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:423" *)
  reg [7:0] vec_data_039_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:424" *)
  reg [7:0] vec_data_039_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:425" *)
  wire [7:0] vec_data_040;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:426" *)
  reg [7:0] vec_data_040_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:427" *)
  reg [7:0] vec_data_040_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:428" *)
  wire [7:0] vec_data_041;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:429" *)
  reg [7:0] vec_data_041_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:430" *)
  reg [7:0] vec_data_041_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:431" *)
  wire [7:0] vec_data_042;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:432" *)
  reg [7:0] vec_data_042_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:433" *)
  reg [7:0] vec_data_042_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:434" *)
  wire [7:0] vec_data_043;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:435" *)
  reg [7:0] vec_data_043_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:436" *)
  reg [7:0] vec_data_043_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:437" *)
  wire [7:0] vec_data_044;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:438" *)
  reg [7:0] vec_data_044_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:439" *)
  reg [7:0] vec_data_044_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:440" *)
  wire [7:0] vec_data_045;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:441" *)
  reg [7:0] vec_data_045_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:442" *)
  reg [7:0] vec_data_045_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:443" *)
  wire [7:0] vec_data_046;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:444" *)
  reg [7:0] vec_data_046_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:445" *)
  reg [7:0] vec_data_046_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:446" *)
  wire [7:0] vec_data_047;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:447" *)
  reg [7:0] vec_data_047_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:448" *)
  reg [7:0] vec_data_047_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:449" *)
  wire [7:0] vec_data_048;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:450" *)
  reg [7:0] vec_data_048_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:451" *)
  reg [7:0] vec_data_048_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:452" *)
  wire [7:0] vec_data_049;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:453" *)
  reg [7:0] vec_data_049_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:454" *)
  reg [7:0] vec_data_049_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:455" *)
  wire [7:0] vec_data_050;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:456" *)
  reg [7:0] vec_data_050_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:457" *)
  reg [7:0] vec_data_050_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:458" *)
  wire [7:0] vec_data_051;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:459" *)
  reg [7:0] vec_data_051_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:460" *)
  reg [7:0] vec_data_051_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:461" *)
  wire [7:0] vec_data_052;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:462" *)
  reg [7:0] vec_data_052_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:463" *)
  reg [7:0] vec_data_052_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:464" *)
  wire [7:0] vec_data_053;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:465" *)
  reg [7:0] vec_data_053_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:466" *)
  reg [7:0] vec_data_053_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:467" *)
  wire [7:0] vec_data_054;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:468" *)
  reg [7:0] vec_data_054_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:469" *)
  reg [7:0] vec_data_054_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:470" *)
  wire [7:0] vec_data_055;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:471" *)
  reg [7:0] vec_data_055_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:472" *)
  reg [7:0] vec_data_055_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:473" *)
  wire [7:0] vec_data_056;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:474" *)
  reg [7:0] vec_data_056_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:475" *)
  reg [7:0] vec_data_056_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:476" *)
  wire [7:0] vec_data_057;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:477" *)
  reg [7:0] vec_data_057_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:478" *)
  reg [7:0] vec_data_057_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:479" *)
  wire [7:0] vec_data_058;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:480" *)
  reg [7:0] vec_data_058_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:481" *)
  reg [7:0] vec_data_058_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:482" *)
  wire [7:0] vec_data_059;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:483" *)
  reg [7:0] vec_data_059_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:484" *)
  reg [7:0] vec_data_059_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:485" *)
  wire [7:0] vec_data_060;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:486" *)
  reg [7:0] vec_data_060_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:487" *)
  reg [7:0] vec_data_060_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:488" *)
  wire [7:0] vec_data_061;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:489" *)
  reg [7:0] vec_data_061_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:490" *)
  reg [7:0] vec_data_061_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:491" *)
  wire [7:0] vec_data_062;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:492" *)
  reg [7:0] vec_data_062_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:493" *)
  reg [7:0] vec_data_062_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:494" *)
  wire [7:0] vec_data_063;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:495" *)
  reg [7:0] vec_data_063_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:496" *)
  reg [7:0] vec_data_063_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:497" *)
  wire [7:0] vec_data_064;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:498" *)
  reg [7:0] vec_data_064_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:499" *)
  reg [7:0] vec_data_064_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:500" *)
  wire [7:0] vec_data_065;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:501" *)
  reg [7:0] vec_data_065_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:502" *)
  reg [7:0] vec_data_065_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:503" *)
  wire [7:0] vec_data_066;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:504" *)
  reg [7:0] vec_data_066_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:505" *)
  reg [7:0] vec_data_066_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:506" *)
  wire [7:0] vec_data_067;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:507" *)
  reg [7:0] vec_data_067_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:508" *)
  reg [7:0] vec_data_067_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:509" *)
  wire [7:0] vec_data_068;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:510" *)
  reg [7:0] vec_data_068_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:511" *)
  reg [7:0] vec_data_068_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:512" *)
  wire [7:0] vec_data_069;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:513" *)
  reg [7:0] vec_data_069_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:514" *)
  reg [7:0] vec_data_069_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:515" *)
  wire [7:0] vec_data_070;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:516" *)
  reg [7:0] vec_data_070_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:517" *)
  reg [7:0] vec_data_070_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:518" *)
  wire [7:0] vec_data_071;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:519" *)
  reg [7:0] vec_data_071_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:520" *)
  reg [7:0] vec_data_071_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:521" *)
  wire [7:0] vec_data_072;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:522" *)
  reg [7:0] vec_data_072_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:523" *)
  reg [7:0] vec_data_072_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:524" *)
  wire [7:0] vec_data_073;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:525" *)
  reg [7:0] vec_data_073_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:526" *)
  reg [7:0] vec_data_073_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:527" *)
  wire [7:0] vec_data_074;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:528" *)
  reg [7:0] vec_data_074_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:529" *)
  reg [7:0] vec_data_074_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:530" *)
  wire [7:0] vec_data_075;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:531" *)
  reg [7:0] vec_data_075_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:532" *)
  reg [7:0] vec_data_075_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:533" *)
  wire [7:0] vec_data_076;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:534" *)
  reg [7:0] vec_data_076_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:535" *)
  reg [7:0] vec_data_076_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:536" *)
  wire [7:0] vec_data_077;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:537" *)
  reg [7:0] vec_data_077_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:538" *)
  reg [7:0] vec_data_077_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:539" *)
  wire [7:0] vec_data_078;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:540" *)
  reg [7:0] vec_data_078_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:541" *)
  reg [7:0] vec_data_078_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:542" *)
  wire [7:0] vec_data_079;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:543" *)
  reg [7:0] vec_data_079_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:544" *)
  reg [7:0] vec_data_079_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:545" *)
  wire [7:0] vec_data_080;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:546" *)
  reg [7:0] vec_data_080_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:547" *)
  reg [7:0] vec_data_080_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:548" *)
  wire [7:0] vec_data_081;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:549" *)
  reg [7:0] vec_data_081_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:550" *)
  reg [7:0] vec_data_081_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:551" *)
  wire [7:0] vec_data_082;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:552" *)
  reg [7:0] vec_data_082_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:553" *)
  reg [7:0] vec_data_082_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:554" *)
  wire [7:0] vec_data_083;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:555" *)
  reg [7:0] vec_data_083_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:556" *)
  reg [7:0] vec_data_083_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:557" *)
  wire [7:0] vec_data_084;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:558" *)
  reg [7:0] vec_data_084_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:559" *)
  reg [7:0] vec_data_084_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:560" *)
  wire [7:0] vec_data_085;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:561" *)
  reg [7:0] vec_data_085_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:562" *)
  reg [7:0] vec_data_085_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:563" *)
  wire [7:0] vec_data_086;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:564" *)
  reg [7:0] vec_data_086_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:565" *)
  reg [7:0] vec_data_086_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:566" *)
  wire [7:0] vec_data_087;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:567" *)
  reg [7:0] vec_data_087_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:568" *)
  reg [7:0] vec_data_087_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:569" *)
  wire [7:0] vec_data_088;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:570" *)
  reg [7:0] vec_data_088_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:571" *)
  reg [7:0] vec_data_088_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:572" *)
  wire [7:0] vec_data_089;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:573" *)
  reg [7:0] vec_data_089_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:574" *)
  reg [7:0] vec_data_089_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:575" *)
  wire [7:0] vec_data_090;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:576" *)
  reg [7:0] vec_data_090_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:577" *)
  reg [7:0] vec_data_090_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:578" *)
  wire [7:0] vec_data_091;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:579" *)
  reg [7:0] vec_data_091_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:580" *)
  reg [7:0] vec_data_091_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:581" *)
  wire [7:0] vec_data_092;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:582" *)
  reg [7:0] vec_data_092_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:583" *)
  reg [7:0] vec_data_092_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:584" *)
  wire [7:0] vec_data_093;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:585" *)
  reg [7:0] vec_data_093_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:586" *)
  reg [7:0] vec_data_093_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:587" *)
  wire [7:0] vec_data_094;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:588" *)
  reg [7:0] vec_data_094_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:589" *)
  reg [7:0] vec_data_094_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:590" *)
  wire [7:0] vec_data_095;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:591" *)
  reg [7:0] vec_data_095_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:592" *)
  reg [7:0] vec_data_095_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:593" *)
  wire [7:0] vec_data_096;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:594" *)
  reg [7:0] vec_data_096_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:595" *)
  reg [7:0] vec_data_096_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:596" *)
  wire [7:0] vec_data_097;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:597" *)
  reg [7:0] vec_data_097_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:598" *)
  reg [7:0] vec_data_097_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:599" *)
  wire [7:0] vec_data_098;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:600" *)
  reg [7:0] vec_data_098_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:601" *)
  reg [7:0] vec_data_098_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:602" *)
  wire [7:0] vec_data_099;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:603" *)
  reg [7:0] vec_data_099_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:604" *)
  reg [7:0] vec_data_099_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:605" *)
  wire [7:0] vec_data_100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:606" *)
  reg [7:0] vec_data_100_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:607" *)
  reg [7:0] vec_data_100_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:608" *)
  wire [7:0] vec_data_101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:609" *)
  reg [7:0] vec_data_101_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:610" *)
  reg [7:0] vec_data_101_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:611" *)
  wire [7:0] vec_data_102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:612" *)
  reg [7:0] vec_data_102_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:613" *)
  reg [7:0] vec_data_102_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:614" *)
  wire [7:0] vec_data_103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:615" *)
  reg [7:0] vec_data_103_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:616" *)
  reg [7:0] vec_data_103_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:617" *)
  wire [7:0] vec_data_104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:618" *)
  reg [7:0] vec_data_104_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:619" *)
  reg [7:0] vec_data_104_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:620" *)
  wire [7:0] vec_data_105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:621" *)
  reg [7:0] vec_data_105_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:622" *)
  reg [7:0] vec_data_105_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:623" *)
  wire [7:0] vec_data_106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:624" *)
  reg [7:0] vec_data_106_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:625" *)
  reg [7:0] vec_data_106_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:626" *)
  wire [7:0] vec_data_107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:627" *)
  reg [7:0] vec_data_107_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:628" *)
  reg [7:0] vec_data_107_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:629" *)
  wire [7:0] vec_data_108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:630" *)
  reg [7:0] vec_data_108_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:631" *)
  reg [7:0] vec_data_108_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:632" *)
  wire [7:0] vec_data_109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:633" *)
  reg [7:0] vec_data_109_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:634" *)
  reg [7:0] vec_data_109_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:635" *)
  wire [7:0] vec_data_110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:636" *)
  reg [7:0] vec_data_110_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:637" *)
  reg [7:0] vec_data_110_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:638" *)
  wire [7:0] vec_data_111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:639" *)
  reg [7:0] vec_data_111_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:640" *)
  reg [7:0] vec_data_111_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:641" *)
  wire [7:0] vec_data_112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:642" *)
  reg [7:0] vec_data_112_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:643" *)
  reg [7:0] vec_data_112_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:644" *)
  wire [7:0] vec_data_113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:645" *)
  reg [7:0] vec_data_113_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:646" *)
  reg [7:0] vec_data_113_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:647" *)
  wire [7:0] vec_data_114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:648" *)
  reg [7:0] vec_data_114_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:649" *)
  reg [7:0] vec_data_114_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:650" *)
  wire [7:0] vec_data_115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:651" *)
  reg [7:0] vec_data_115_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:652" *)
  reg [7:0] vec_data_115_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:653" *)
  wire [7:0] vec_data_116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:654" *)
  reg [7:0] vec_data_116_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:655" *)
  reg [7:0] vec_data_116_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:656" *)
  wire [7:0] vec_data_117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:657" *)
  reg [7:0] vec_data_117_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:658" *)
  reg [7:0] vec_data_117_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:659" *)
  wire [7:0] vec_data_118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:660" *)
  reg [7:0] vec_data_118_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:661" *)
  reg [7:0] vec_data_118_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:662" *)
  wire [7:0] vec_data_119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:663" *)
  reg [7:0] vec_data_119_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:664" *)
  reg [7:0] vec_data_119_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:665" *)
  wire [7:0] vec_data_120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:666" *)
  reg [7:0] vec_data_120_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:667" *)
  reg [7:0] vec_data_120_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:668" *)
  wire [7:0] vec_data_121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:669" *)
  reg [7:0] vec_data_121_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:670" *)
  reg [7:0] vec_data_121_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:671" *)
  wire [7:0] vec_data_122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:672" *)
  reg [7:0] vec_data_122_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:673" *)
  reg [7:0] vec_data_122_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:674" *)
  wire [7:0] vec_data_123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:675" *)
  reg [7:0] vec_data_123_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:676" *)
  reg [7:0] vec_data_123_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:677" *)
  wire [7:0] vec_data_124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:678" *)
  reg [7:0] vec_data_124_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:679" *)
  reg [7:0] vec_data_124_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:680" *)
  wire [7:0] vec_data_125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:681" *)
  reg [7:0] vec_data_125_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:682" *)
  reg [7:0] vec_data_125_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:683" *)
  wire [7:0] vec_data_126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:684" *)
  reg [7:0] vec_data_126_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:685" *)
  reg [7:0] vec_data_126_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:686" *)
  wire [7:0] vec_data_127;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:687" *)
  reg [7:0] vec_data_127_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:688" *)
  reg [7:0] vec_data_127_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:689" *)
  wire vec_sum_000;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:690" *)
  reg vec_sum_000_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:691" *)
  wire [1:0] vec_sum_001;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:692" *)
  reg [1:0] vec_sum_001_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:693" *)
  wire [1:0] vec_sum_002;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:694" *)
  reg [1:0] vec_sum_002_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:695" *)
  wire [2:0] vec_sum_003;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:696" *)
  reg [2:0] vec_sum_003_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:697" *)
  wire [2:0] vec_sum_004;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:698" *)
  reg [2:0] vec_sum_004_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:699" *)
  wire [2:0] vec_sum_005;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:700" *)
  reg [2:0] vec_sum_005_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:701" *)
  wire [2:0] vec_sum_006;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:702" *)
  reg [2:0] vec_sum_006_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:703" *)
  wire [3:0] vec_sum_007;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:704" *)
  reg [3:0] vec_sum_007_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:705" *)
  wire [3:0] vec_sum_008;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:706" *)
  reg [3:0] vec_sum_008_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:707" *)
  wire [3:0] vec_sum_009;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:708" *)
  reg [3:0] vec_sum_009_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:709" *)
  wire [3:0] vec_sum_010;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:710" *)
  reg [3:0] vec_sum_010_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:711" *)
  wire [3:0] vec_sum_011;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:712" *)
  reg [3:0] vec_sum_011_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:713" *)
  wire [3:0] vec_sum_012;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:714" *)
  reg [3:0] vec_sum_012_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:715" *)
  wire [3:0] vec_sum_013;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:716" *)
  reg [3:0] vec_sum_013_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:717" *)
  wire [3:0] vec_sum_014;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:718" *)
  reg [3:0] vec_sum_014_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:719" *)
  wire [4:0] vec_sum_015;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:720" *)
  reg [4:0] vec_sum_015_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:721" *)
  wire [4:0] vec_sum_016;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:722" *)
  reg [4:0] vec_sum_016_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:723" *)
  wire [4:0] vec_sum_017;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:724" *)
  reg [4:0] vec_sum_017_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:725" *)
  wire [4:0] vec_sum_018;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:726" *)
  reg [4:0] vec_sum_018_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:727" *)
  wire [4:0] vec_sum_019;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:728" *)
  reg [4:0] vec_sum_019_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:729" *)
  wire [4:0] vec_sum_020;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:730" *)
  reg [4:0] vec_sum_020_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:731" *)
  wire [4:0] vec_sum_021;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:732" *)
  reg [4:0] vec_sum_021_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:733" *)
  wire [4:0] vec_sum_022;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:734" *)
  reg [4:0] vec_sum_022_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:735" *)
  wire [4:0] vec_sum_023;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:736" *)
  reg [4:0] vec_sum_023_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:737" *)
  wire [4:0] vec_sum_024;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:738" *)
  reg [4:0] vec_sum_024_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:739" *)
  wire [4:0] vec_sum_025;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:740" *)
  reg [4:0] vec_sum_025_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:741" *)
  wire [4:0] vec_sum_026;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:742" *)
  reg [4:0] vec_sum_026_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:743" *)
  wire [4:0] vec_sum_027;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:744" *)
  reg [4:0] vec_sum_027_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:745" *)
  wire [4:0] vec_sum_028;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:746" *)
  reg [4:0] vec_sum_028_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:747" *)
  wire [4:0] vec_sum_029;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:748" *)
  reg [4:0] vec_sum_029_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:749" *)
  wire [4:0] vec_sum_030;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:750" *)
  reg [4:0] vec_sum_030_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:751" *)
  wire [5:0] vec_sum_031;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:752" *)
  reg [5:0] vec_sum_031_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:753" *)
  wire [5:0] vec_sum_032;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:754" *)
  reg [5:0] vec_sum_032_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:755" *)
  wire [5:0] vec_sum_033;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:756" *)
  reg [5:0] vec_sum_033_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:757" *)
  wire [5:0] vec_sum_034;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:758" *)
  reg [5:0] vec_sum_034_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:759" *)
  wire [5:0] vec_sum_035;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:760" *)
  reg [5:0] vec_sum_035_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:761" *)
  wire [5:0] vec_sum_036;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:762" *)
  reg [5:0] vec_sum_036_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:763" *)
  wire [5:0] vec_sum_037;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:764" *)
  reg [5:0] vec_sum_037_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:765" *)
  wire [5:0] vec_sum_038;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:766" *)
  reg [5:0] vec_sum_038_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:767" *)
  wire [5:0] vec_sum_039;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:768" *)
  reg [5:0] vec_sum_039_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:769" *)
  wire [5:0] vec_sum_040;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:770" *)
  reg [5:0] vec_sum_040_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:771" *)
  wire [5:0] vec_sum_041;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:772" *)
  reg [5:0] vec_sum_041_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:773" *)
  wire [5:0] vec_sum_042;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:774" *)
  reg [5:0] vec_sum_042_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:775" *)
  wire [5:0] vec_sum_043;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:776" *)
  reg [5:0] vec_sum_043_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:777" *)
  wire [5:0] vec_sum_044;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:778" *)
  reg [5:0] vec_sum_044_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:779" *)
  wire [5:0] vec_sum_045;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:780" *)
  reg [5:0] vec_sum_045_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:781" *)
  wire [5:0] vec_sum_046;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:782" *)
  reg [5:0] vec_sum_046_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:783" *)
  wire [5:0] vec_sum_047;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:784" *)
  reg [5:0] vec_sum_047_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:785" *)
  wire [5:0] vec_sum_048;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:786" *)
  reg [5:0] vec_sum_048_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:787" *)
  wire [5:0] vec_sum_049;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:788" *)
  reg [5:0] vec_sum_049_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:789" *)
  wire [5:0] vec_sum_050;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:790" *)
  reg [5:0] vec_sum_050_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:791" *)
  wire [5:0] vec_sum_051;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:792" *)
  reg [5:0] vec_sum_051_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:793" *)
  wire [5:0] vec_sum_052;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:794" *)
  reg [5:0] vec_sum_052_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:795" *)
  wire [5:0] vec_sum_053;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:796" *)
  reg [5:0] vec_sum_053_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:797" *)
  wire [5:0] vec_sum_054;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:798" *)
  reg [5:0] vec_sum_054_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:799" *)
  wire [5:0] vec_sum_055;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:800" *)
  reg [5:0] vec_sum_055_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:801" *)
  wire [5:0] vec_sum_056;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:802" *)
  reg [5:0] vec_sum_056_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:803" *)
  wire [5:0] vec_sum_057;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:804" *)
  reg [5:0] vec_sum_057_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:805" *)
  wire [5:0] vec_sum_058;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:806" *)
  reg [5:0] vec_sum_058_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:807" *)
  wire [5:0] vec_sum_059;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:808" *)
  reg [5:0] vec_sum_059_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:809" *)
  wire [5:0] vec_sum_060;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:810" *)
  reg [5:0] vec_sum_060_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:811" *)
  wire [5:0] vec_sum_061;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:812" *)
  reg [5:0] vec_sum_061_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:813" *)
  wire [5:0] vec_sum_062;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:814" *)
  reg [5:0] vec_sum_062_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:815" *)
  wire [6:0] vec_sum_063;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:816" *)
  reg [6:0] vec_sum_063_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:817" *)
  wire [6:0] vec_sum_064;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:818" *)
  reg [6:0] vec_sum_064_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:819" *)
  wire [6:0] vec_sum_065;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:820" *)
  reg [6:0] vec_sum_065_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:821" *)
  wire [6:0] vec_sum_066;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:822" *)
  reg [6:0] vec_sum_066_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:823" *)
  wire [6:0] vec_sum_067;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:824" *)
  reg [6:0] vec_sum_067_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:825" *)
  wire [6:0] vec_sum_068;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:826" *)
  reg [6:0] vec_sum_068_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:827" *)
  wire [6:0] vec_sum_069;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:828" *)
  reg [6:0] vec_sum_069_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:829" *)
  wire [6:0] vec_sum_070;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:830" *)
  reg [6:0] vec_sum_070_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:831" *)
  wire [6:0] vec_sum_071;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:832" *)
  reg [6:0] vec_sum_071_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:833" *)
  wire [6:0] vec_sum_072;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:834" *)
  reg [6:0] vec_sum_072_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:835" *)
  wire [6:0] vec_sum_073;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:836" *)
  reg [6:0] vec_sum_073_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:837" *)
  wire [6:0] vec_sum_074;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:838" *)
  reg [6:0] vec_sum_074_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:839" *)
  wire [6:0] vec_sum_075;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:840" *)
  reg [6:0] vec_sum_075_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:841" *)
  wire [6:0] vec_sum_076;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:842" *)
  reg [6:0] vec_sum_076_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:843" *)
  wire [6:0] vec_sum_077;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:844" *)
  reg [6:0] vec_sum_077_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:845" *)
  wire [6:0] vec_sum_078;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:846" *)
  reg [6:0] vec_sum_078_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:847" *)
  wire [6:0] vec_sum_079;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:848" *)
  reg [6:0] vec_sum_079_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:849" *)
  wire [6:0] vec_sum_080;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:850" *)
  reg [6:0] vec_sum_080_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:851" *)
  wire [6:0] vec_sum_081;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:852" *)
  reg [6:0] vec_sum_081_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:853" *)
  wire [6:0] vec_sum_082;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:854" *)
  reg [6:0] vec_sum_082_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:855" *)
  wire [6:0] vec_sum_083;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:856" *)
  reg [6:0] vec_sum_083_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:857" *)
  wire [6:0] vec_sum_084;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:858" *)
  reg [6:0] vec_sum_084_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:859" *)
  wire [6:0] vec_sum_085;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:860" *)
  reg [6:0] vec_sum_085_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:861" *)
  wire [6:0] vec_sum_086;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:862" *)
  reg [6:0] vec_sum_086_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:863" *)
  wire [6:0] vec_sum_087;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:864" *)
  reg [6:0] vec_sum_087_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:865" *)
  wire [6:0] vec_sum_088;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:866" *)
  reg [6:0] vec_sum_088_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:867" *)
  wire [6:0] vec_sum_089;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:868" *)
  reg [6:0] vec_sum_089_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:869" *)
  wire [6:0] vec_sum_090;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:870" *)
  reg [6:0] vec_sum_090_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:871" *)
  wire [6:0] vec_sum_091;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:872" *)
  reg [6:0] vec_sum_091_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:873" *)
  wire [6:0] vec_sum_092;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:874" *)
  reg [6:0] vec_sum_092_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:875" *)
  wire [6:0] vec_sum_093;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:876" *)
  reg [6:0] vec_sum_093_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:877" *)
  wire [6:0] vec_sum_094;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:878" *)
  reg [6:0] vec_sum_094_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:879" *)
  wire [6:0] vec_sum_095;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:880" *)
  reg [6:0] vec_sum_095_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:881" *)
  wire [6:0] vec_sum_096;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:882" *)
  reg [6:0] vec_sum_096_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:883" *)
  wire [6:0] vec_sum_097;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:884" *)
  reg [6:0] vec_sum_097_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:885" *)
  wire [6:0] vec_sum_098;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:886" *)
  reg [6:0] vec_sum_098_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:887" *)
  wire [6:0] vec_sum_099;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:888" *)
  reg [6:0] vec_sum_099_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:889" *)
  wire [6:0] vec_sum_100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:890" *)
  reg [6:0] vec_sum_100_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:891" *)
  wire [6:0] vec_sum_101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:892" *)
  reg [6:0] vec_sum_101_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:893" *)
  wire [6:0] vec_sum_102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:894" *)
  reg [6:0] vec_sum_102_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:895" *)
  wire [6:0] vec_sum_103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:896" *)
  reg [6:0] vec_sum_103_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:897" *)
  wire [6:0] vec_sum_104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:898" *)
  reg [6:0] vec_sum_104_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:899" *)
  wire [6:0] vec_sum_105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:900" *)
  reg [6:0] vec_sum_105_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:901" *)
  wire [6:0] vec_sum_106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:902" *)
  reg [6:0] vec_sum_106_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:903" *)
  wire [6:0] vec_sum_107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:904" *)
  reg [6:0] vec_sum_107_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:905" *)
  wire [6:0] vec_sum_108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:906" *)
  reg [6:0] vec_sum_108_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:907" *)
  wire [6:0] vec_sum_109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:908" *)
  reg [6:0] vec_sum_109_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:909" *)
  wire [6:0] vec_sum_110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:910" *)
  reg [6:0] vec_sum_110_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:911" *)
  wire [6:0] vec_sum_111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:912" *)
  reg [6:0] vec_sum_111_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:913" *)
  wire [6:0] vec_sum_112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:914" *)
  reg [6:0] vec_sum_112_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:915" *)
  wire [6:0] vec_sum_113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:916" *)
  reg [6:0] vec_sum_113_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:917" *)
  wire [6:0] vec_sum_114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:918" *)
  reg [6:0] vec_sum_114_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:919" *)
  wire [6:0] vec_sum_115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:920" *)
  reg [6:0] vec_sum_115_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:921" *)
  wire [6:0] vec_sum_116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:922" *)
  reg [6:0] vec_sum_116_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:923" *)
  wire [6:0] vec_sum_117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:924" *)
  reg [6:0] vec_sum_117_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:925" *)
  wire [6:0] vec_sum_118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:926" *)
  reg [6:0] vec_sum_118_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:927" *)
  wire [6:0] vec_sum_119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:928" *)
  reg [6:0] vec_sum_119_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:929" *)
  wire [6:0] vec_sum_120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:930" *)
  reg [6:0] vec_sum_120_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:931" *)
  wire [6:0] vec_sum_121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:932" *)
  reg [6:0] vec_sum_121_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:933" *)
  wire [6:0] vec_sum_122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:934" *)
  reg [6:0] vec_sum_122_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:935" *)
  wire [6:0] vec_sum_123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:936" *)
  reg [6:0] vec_sum_123_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:937" *)
  wire [6:0] vec_sum_124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:938" *)
  reg [6:0] vec_sum_124_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:939" *)
  wire [6:0] vec_sum_125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:940" *)
  reg [6:0] vec_sum_125_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:941" *)
  wire [6:0] vec_sum_126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:942" *)
  reg [6:0] vec_sum_126_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:943" *)
  wire [7:0] vec_sum_127;
  wire [6:0] vec_sum_127_d1;
  assign vec_sum_001 = input_mask_gated[0] + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[1];
  assign _00390_ = vec_sum_001 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[2];
  assign vec_sum_003 = _00390_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[3];
  assign vec_sum_004 = vec_sum_003 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[4];
  assign vec_sum_005 = vec_sum_004 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[5];
  assign vec_sum_006 = vec_sum_005 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1000" *) input_mask_gated[6];
  assign _00391_ = _00390_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *) input_mask_gated[3];
  assign _00392_ = _00391_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *) input_mask_gated[4];
  assign _00393_ = _00392_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *) input_mask_gated[5];
  assign _00394_ = _00393_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *) input_mask_gated[6];
  assign vec_sum_007 = _00394_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1005" *) input_mask_gated[7];
  assign vec_sum_008 = vec_sum_007 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1011" *) input_mask_gated[8];
  assign vec_sum_009 = vec_sum_008 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1017" *) input_mask_gated[9];
  assign vec_sum_010 = vec_sum_009 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1023" *) input_mask_gated[10];
  assign vec_sum_011 = vec_sum_010 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1029" *) input_mask_gated[11];
  assign vec_sum_012 = vec_sum_011 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1035" *) input_mask_gated[12];
  assign vec_sum_013 = vec_sum_012 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1041" *) input_mask_gated[13];
  assign vec_sum_014 = vec_sum_013 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1047" *) input_mask_gated[14];
  assign _00395_ = _00391_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *) input_mask_gated[4];
  assign _00396_ = _00395_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *) input_mask_gated[5];
  assign _00397_ = _00396_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1052" *) input_mask_gated[6];
  assign _00398_ = _00397_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[7];
  assign _00399_ = _00398_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[8];
  assign _00400_ = _00399_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[9];
  assign _00401_ = _00400_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[10];
  assign _00402_ = _00401_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[11];
  assign _00403_ = _00402_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[12];
  assign _00404_ = _00403_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[13];
  assign _00405_ = _00404_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[14];
  assign vec_sum_015 = _00405_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1053" *) input_mask_gated[15];
  assign vec_sum_016 = vec_sum_015 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1060" *) input_mask_gated[16];
  assign vec_sum_017 = vec_sum_016 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1067" *) input_mask_gated[17];
  assign vec_sum_018 = vec_sum_017 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1074" *) input_mask_gated[18];
  assign vec_sum_019 = vec_sum_018 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1081" *) input_mask_gated[19];
  assign vec_sum_020 = vec_sum_019 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1088" *) input_mask_gated[20];
  assign vec_sum_021 = vec_sum_020 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1095" *) input_mask_gated[21];
  assign vec_sum_022 = vec_sum_021 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1102" *) input_mask_gated[22];
  assign vec_sum_023 = vec_sum_022 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1109" *) input_mask_gated[23];
  assign vec_sum_024 = vec_sum_023 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1117" *) input_mask_gated[24];
  assign vec_sum_025 = vec_sum_024 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1125" *) input_mask_gated[25];
  assign vec_sum_026 = vec_sum_025 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1133" *) input_mask_gated[26];
  assign vec_sum_027 = vec_sum_026 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1141" *) input_mask_gated[27];
  assign vec_sum_028 = vec_sum_027 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1149" *) input_mask_gated[28];
  assign vec_sum_029 = vec_sum_028 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1157" *) input_mask_gated[29];
  assign vec_sum_030 = vec_sum_029 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1165" *) input_mask_gated[30];
  assign _00406_ = _00395_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1170" *) input_mask_gated[5];
  assign _00407_ = _00406_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1170" *) input_mask_gated[6];
  assign _00408_ = _00407_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[7];
  assign _00409_ = _00408_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[8];
  assign _00410_ = _00409_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[9];
  assign _00411_ = _00410_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[10];
  assign _00412_ = _00411_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[11];
  assign _00413_ = _00412_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[12];
  assign _00414_ = _00413_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[13];
  assign _00415_ = _00414_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1171" *) input_mask_gated[14];
  assign _00416_ = _00415_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[15];
  assign _00417_ = _00416_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[16];
  assign _00418_ = _00417_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[17];
  assign _00419_ = _00418_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[18];
  assign _00420_ = _00419_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[19];
  assign _00421_ = _00420_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[20];
  assign _00422_ = _00421_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[21];
  assign _00423_ = _00422_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1172" *) input_mask_gated[22];
  assign _00424_ = _00423_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[23];
  assign _00425_ = _00424_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[24];
  assign _00426_ = _00425_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[25];
  assign _00427_ = _00426_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[26];
  assign _00428_ = _00427_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[27];
  assign _00429_ = _00428_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[28];
  assign _00430_ = _00429_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[29];
  assign _00431_ = _00430_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[30];
  assign vec_sum_031 = _00431_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1173" *) input_mask_gated[31];
  assign vec_sum_032 = vec_sum_031 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1182" *) input_mask_gated[32];
  assign vec_sum_033 = vec_sum_032 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1191" *) input_mask_gated[33];
  assign vec_sum_034 = vec_sum_033 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1200" *) input_mask_gated[34];
  assign vec_sum_035 = vec_sum_034 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1209" *) input_mask_gated[35];
  assign vec_sum_036 = vec_sum_035 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1218" *) input_mask_gated[36];
  assign vec_sum_037 = vec_sum_036 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1227" *) input_mask_gated[37];
  assign vec_sum_038 = vec_sum_037 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1236" *) input_mask_gated[38];
  assign vec_sum_039 = vec_sum_038 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1245" *) input_mask_gated[39];
  assign vec_sum_040 = vec_sum_039 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1255" *) input_mask_gated[40];
  assign vec_sum_041 = vec_sum_040 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1265" *) input_mask_gated[41];
  assign vec_sum_042 = vec_sum_041 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1275" *) input_mask_gated[42];
  assign vec_sum_043 = vec_sum_042 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1285" *) input_mask_gated[43];
  assign vec_sum_044 = vec_sum_043 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1295" *) input_mask_gated[44];
  assign vec_sum_045 = vec_sum_044 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1305" *) input_mask_gated[45];
  assign vec_sum_046 = vec_sum_045 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1315" *) input_mask_gated[46];
  assign vec_sum_047 = vec_sum_046 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1325" *) input_mask_gated[47];
  assign vec_sum_048 = vec_sum_047 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1336" *) input_mask_gated[48];
  assign vec_sum_049 = vec_sum_048 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1347" *) input_mask_gated[49];
  assign vec_sum_050 = vec_sum_049 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1358" *) input_mask_gated[50];
  assign vec_sum_051 = vec_sum_050 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1369" *) input_mask_gated[51];
  assign vec_sum_052 = vec_sum_051 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1380" *) input_mask_gated[52];
  assign vec_sum_053 = vec_sum_052 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1391" *) input_mask_gated[53];
  assign vec_sum_054 = vec_sum_053 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1402" *) input_mask_gated[54];
  assign vec_sum_055 = vec_sum_054 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1413" *) input_mask_gated[55];
  assign vec_sum_056 = vec_sum_055 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1425" *) input_mask_gated[56];
  assign vec_sum_057 = vec_sum_056 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1437" *) input_mask_gated[57];
  assign vec_sum_058 = vec_sum_057 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1449" *) input_mask_gated[58];
  assign vec_sum_059 = vec_sum_058 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1461" *) input_mask_gated[59];
  assign vec_sum_060 = vec_sum_059 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1473" *) input_mask_gated[60];
  assign vec_sum_061 = vec_sum_060 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1485" *) input_mask_gated[61];
  assign vec_sum_062 = vec_sum_061 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1497" *) input_mask_gated[62];
  assign _00432_ = _00406_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1502" *) input_mask_gated[6];
  assign _00433_ = _00432_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[7];
  assign _00434_ = _00433_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[8];
  assign _00435_ = _00434_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[9];
  assign _00436_ = _00435_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[10];
  assign _00437_ = _00436_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[11];
  assign _00438_ = _00437_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[12];
  assign _00439_ = _00438_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[13];
  assign _00440_ = _00439_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1503" *) input_mask_gated[14];
  assign _00441_ = _00440_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[15];
  assign _00442_ = _00441_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[16];
  assign _00443_ = _00442_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[17];
  assign _00444_ = _00443_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[18];
  assign _00445_ = _00444_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[19];
  assign _00446_ = _00445_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[20];
  assign _00447_ = _00446_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[21];
  assign _00448_ = _00447_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1504" *) input_mask_gated[22];
  assign _00449_ = _00448_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[23];
  assign _00450_ = _00449_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[24];
  assign _00451_ = _00450_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[25];
  assign _00452_ = _00451_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[26];
  assign _00453_ = _00452_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[27];
  assign _00454_ = _00453_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[28];
  assign _00455_ = _00454_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[29];
  assign _00456_ = _00455_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1505" *) input_mask_gated[30];
  assign _00457_ = _00456_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[31];
  assign _00458_ = _00457_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[32];
  assign _00459_ = _00458_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[33];
  assign _00460_ = _00459_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[34];
  assign _00461_ = _00460_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[35];
  assign _00462_ = _00461_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[36];
  assign _00463_ = _00462_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[37];
  assign _00464_ = _00463_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1506" *) input_mask_gated[38];
  assign _00465_ = _00464_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[39];
  assign _00466_ = _00465_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[40];
  assign _00467_ = _00466_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[41];
  assign _00468_ = _00467_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[42];
  assign _00469_ = _00468_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[43];
  assign _00470_ = _00469_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[44];
  assign _00471_ = _00470_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[45];
  assign _00472_ = _00471_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1507" *) input_mask_gated[46];
  assign _00473_ = _00472_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[47];
  assign _00474_ = _00473_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[48];
  assign _00475_ = _00474_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[49];
  assign _00476_ = _00475_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[50];
  assign _00477_ = _00476_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[51];
  assign _00478_ = _00477_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[52];
  assign _00479_ = _00478_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[53];
  assign _00480_ = _00479_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1508" *) input_mask_gated[54];
  assign _00481_ = _00480_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[55];
  assign _00482_ = _00481_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[56];
  assign _00483_ = _00482_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[57];
  assign _00484_ = _00483_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[58];
  assign _00485_ = _00484_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[59];
  assign _00486_ = _00485_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[60];
  assign _00487_ = _00486_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[61];
  assign _00488_ = _00487_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[62];
  assign vec_sum_063 = _00488_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1509" *) input_mask_gated[63];
  assign vec_sum_064 = vec_sum_063 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1522" *) input_mask_gated[64];
  assign vec_sum_065 = vec_sum_064 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1535" *) input_mask_gated[65];
  assign vec_sum_066 = vec_sum_065 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1548" *) input_mask_gated[66];
  assign vec_sum_067 = vec_sum_066 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1561" *) input_mask_gated[67];
  assign vec_sum_068 = vec_sum_067 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1574" *) input_mask_gated[68];
  assign vec_sum_069 = vec_sum_068 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1587" *) input_mask_gated[69];
  assign vec_sum_070 = vec_sum_069 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1600" *) input_mask_gated[70];
  assign vec_sum_071 = vec_sum_070 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1613" *) input_mask_gated[71];
  assign vec_sum_072 = vec_sum_071 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1627" *) input_mask_gated[72];
  assign vec_sum_073 = vec_sum_072 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1641" *) input_mask_gated[73];
  assign vec_sum_074 = vec_sum_073 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1655" *) input_mask_gated[74];
  assign vec_sum_075 = vec_sum_074 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1669" *) input_mask_gated[75];
  assign vec_sum_076 = vec_sum_075 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1683" *) input_mask_gated[76];
  assign vec_sum_077 = vec_sum_076 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1697" *) input_mask_gated[77];
  assign vec_sum_078 = vec_sum_077 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1711" *) input_mask_gated[78];
  assign vec_sum_079 = vec_sum_078 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1725" *) input_mask_gated[79];
  assign vec_sum_080 = vec_sum_079 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1740" *) input_mask_gated[80];
  assign vec_sum_081 = vec_sum_080 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1755" *) input_mask_gated[81];
  assign vec_sum_082 = vec_sum_081 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1770" *) input_mask_gated[82];
  assign vec_sum_083 = vec_sum_082 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1785" *) input_mask_gated[83];
  assign vec_sum_084 = vec_sum_083 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1800" *) input_mask_gated[84];
  assign vec_sum_085 = vec_sum_084 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1815" *) input_mask_gated[85];
  assign vec_sum_086 = vec_sum_085 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1830" *) input_mask_gated[86];
  assign vec_sum_087 = vec_sum_086 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1845" *) input_mask_gated[87];
  assign vec_sum_088 = vec_sum_087 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1861" *) input_mask_gated[88];
  assign vec_sum_089 = vec_sum_088 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1877" *) input_mask_gated[89];
  assign vec_sum_090 = vec_sum_089 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1893" *) input_mask_gated[90];
  assign vec_sum_091 = vec_sum_090 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1909" *) input_mask_gated[91];
  assign vec_sum_092 = vec_sum_091 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1925" *) input_mask_gated[92];
  assign vec_sum_093 = vec_sum_092 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1941" *) input_mask_gated[93];
  assign vec_sum_094 = vec_sum_093 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1957" *) input_mask_gated[94];
  assign vec_sum_095 = vec_sum_094 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1973" *) input_mask_gated[95];
  assign vec_sum_096 = vec_sum_095 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:1990" *) input_mask_gated[96];
  assign vec_sum_097 = vec_sum_096 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2007" *) input_mask_gated[97];
  assign vec_sum_098 = vec_sum_097 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2024" *) input_mask_gated[98];
  assign vec_sum_099 = vec_sum_098 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2041" *) input_mask_gated[99];
  assign vec_sum_100 = vec_sum_099 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2058" *) input_mask_gated[100];
  assign vec_sum_101 = vec_sum_100 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2075" *) input_mask_gated[101];
  assign vec_sum_102 = vec_sum_101 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2092" *) input_mask_gated[102];
  assign vec_sum_103 = vec_sum_102 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2109" *) input_mask_gated[103];
  assign vec_sum_104 = vec_sum_103 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2127" *) input_mask_gated[104];
  assign vec_sum_105 = vec_sum_104 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2145" *) input_mask_gated[105];
  assign vec_sum_106 = vec_sum_105 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2163" *) input_mask_gated[106];
  assign vec_sum_107 = vec_sum_106 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2181" *) input_mask_gated[107];
  assign vec_sum_108 = vec_sum_107 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2199" *) input_mask_gated[108];
  assign vec_sum_109 = vec_sum_108 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2217" *) input_mask_gated[109];
  assign vec_sum_110 = vec_sum_109 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2235" *) input_mask_gated[110];
  assign vec_sum_111 = vec_sum_110 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2253" *) input_mask_gated[111];
  assign vec_sum_112 = vec_sum_111 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2272" *) input_mask_gated[112];
  assign vec_sum_113 = vec_sum_112 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2291" *) input_mask_gated[113];
  assign vec_sum_114 = vec_sum_113 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2310" *) input_mask_gated[114];
  assign vec_sum_115 = vec_sum_114 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2329" *) input_mask_gated[115];
  assign vec_sum_116 = vec_sum_115 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2348" *) input_mask_gated[116];
  assign vec_sum_117 = vec_sum_116 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2367" *) input_mask_gated[117];
  assign vec_sum_118 = vec_sum_117 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2386" *) input_mask_gated[118];
  assign vec_sum_119 = vec_sum_118 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2405" *) input_mask_gated[119];
  assign vec_sum_120 = vec_sum_119 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2425" *) input_mask_gated[120];
  assign vec_sum_121 = vec_sum_120 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2445" *) input_mask_gated[121];
  assign vec_sum_122 = vec_sum_121 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2465" *) input_mask_gated[122];
  assign vec_sum_123 = vec_sum_122 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2485" *) input_mask_gated[123];
  assign vec_sum_124 = vec_sum_123 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2505" *) input_mask_gated[124];
  assign vec_sum_125 = vec_sum_124 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2525" *) input_mask_gated[125];
  assign vec_sum_126 = vec_sum_125 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2545" *) input_mask_gated[126];
  assign _00489_ = _00432_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[7];
  assign _00490_ = _00489_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[8];
  assign _00491_ = _00490_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[9];
  assign _00492_ = _00491_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[10];
  assign _00493_ = _00492_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[11];
  assign _00494_ = _00493_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[12];
  assign _00495_ = _00494_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[13];
  assign _00496_ = _00495_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2551" *) input_mask_gated[14];
  assign _00497_ = _00496_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[15];
  assign _00498_ = _00497_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[16];
  assign _00499_ = _00498_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[17];
  assign _00500_ = _00499_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[18];
  assign _00501_ = _00500_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[19];
  assign _00502_ = _00501_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[20];
  assign _00503_ = _00502_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[21];
  assign _00504_ = _00503_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2552" *) input_mask_gated[22];
  assign _00505_ = _00504_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[23];
  assign _00506_ = _00505_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[24];
  assign _00507_ = _00506_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[25];
  assign _00508_ = _00507_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[26];
  assign _00509_ = _00508_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[27];
  assign _00510_ = _00509_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[28];
  assign _00511_ = _00510_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[29];
  assign _00512_ = _00511_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2553" *) input_mask_gated[30];
  assign _00513_ = _00512_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[31];
  assign _00514_ = _00513_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[32];
  assign _00515_ = _00514_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[33];
  assign _00516_ = _00515_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[34];
  assign _00517_ = _00516_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[35];
  assign _00518_ = _00517_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[36];
  assign _00519_ = _00518_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[37];
  assign _00520_ = _00519_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2554" *) input_mask_gated[38];
  assign _00521_ = _00520_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[39];
  assign _00522_ = _00521_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[40];
  assign _00523_ = _00522_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[41];
  assign _00524_ = _00523_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[42];
  assign _00525_ = _00524_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[43];
  assign _00526_ = _00525_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[44];
  assign _00527_ = _00526_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[45];
  assign _00528_ = _00527_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2555" *) input_mask_gated[46];
  assign _00529_ = _00528_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[47];
  assign _00530_ = _00529_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[48];
  assign _00531_ = _00530_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[49];
  assign _00532_ = _00531_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[50];
  assign _00533_ = _00532_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[51];
  assign _00534_ = _00533_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[52];
  assign _00535_ = _00534_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[53];
  assign _00536_ = _00535_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2556" *) input_mask_gated[54];
  assign _00537_ = _00536_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[55];
  assign _00538_ = _00537_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[56];
  assign _00539_ = _00538_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[57];
  assign _00540_ = _00539_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[58];
  assign _00541_ = _00540_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[59];
  assign _00542_ = _00541_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[60];
  assign _00543_ = _00542_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[61];
  assign _00544_ = _00543_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2557" *) input_mask_gated[62];
  assign _00545_ = _00544_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[63];
  assign _00546_ = _00545_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[64];
  assign _00547_ = _00546_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[65];
  assign _00548_ = _00547_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[66];
  assign _00549_ = _00548_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[67];
  assign _00550_ = _00549_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[68];
  assign _00551_ = _00550_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[69];
  assign _00552_ = _00551_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2558" *) input_mask_gated[70];
  assign _00553_ = _00552_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[71];
  assign _00554_ = _00553_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[72];
  assign _00555_ = _00554_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[73];
  assign _00556_ = _00555_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[74];
  assign _00557_ = _00556_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[75];
  assign _00558_ = _00557_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[76];
  assign _00559_ = _00558_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[77];
  assign _00560_ = _00559_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2559" *) input_mask_gated[78];
  assign _00561_ = _00560_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[79];
  assign _00562_ = _00561_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[80];
  assign _00563_ = _00562_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[81];
  assign _00564_ = _00563_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[82];
  assign _00565_ = _00564_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[83];
  assign _00566_ = _00565_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[84];
  assign _00567_ = _00566_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[85];
  assign _00568_ = _00567_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2560" *) input_mask_gated[86];
  assign _00569_ = _00568_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[87];
  assign _00570_ = _00569_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[88];
  assign _00571_ = _00570_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[89];
  assign _00572_ = _00571_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[90];
  assign _00573_ = _00572_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[91];
  assign _00574_ = _00573_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[92];
  assign _00575_ = _00574_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[93];
  assign _00576_ = _00575_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2561" *) input_mask_gated[94];
  assign _00577_ = _00576_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[95];
  assign _00578_ = _00577_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[96];
  assign _00579_ = _00578_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[97];
  assign _00580_ = _00579_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[98];
  assign _00581_ = _00580_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[99];
  assign _00582_ = _00581_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[100];
  assign _00583_ = _00582_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[101];
  assign _00584_ = _00583_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2562" *) input_mask_gated[102];
  assign _00585_ = _00584_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[103];
  assign _00586_ = _00585_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[104];
  assign _00587_ = _00586_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[105];
  assign _00588_ = _00587_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[106];
  assign _00589_ = _00588_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[107];
  assign _00590_ = _00589_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[108];
  assign _00591_ = _00590_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[109];
  assign _00592_ = _00591_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2563" *) input_mask_gated[110];
  assign _00593_ = _00592_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[111];
  assign _00594_ = _00593_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[112];
  assign _00595_ = _00594_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[113];
  assign _00596_ = _00595_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[114];
  assign _00597_ = _00596_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[115];
  assign _00598_ = _00597_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[116];
  assign _00599_ = _00598_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[117];
  assign _00600_ = _00599_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2564" *) input_mask_gated[118];
  assign _00601_ = _00600_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[119];
  assign _00602_ = _00601_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[120];
  assign _00603_ = _00602_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[121];
  assign _00604_ = _00603_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[122];
  assign _00605_ = _00604_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[123];
  assign _00606_ = _00605_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[124];
  assign _00607_ = _00606_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[125];
  assign _00608_ = _00607_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[126];
  assign vec_sum_127 = _00608_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2565" *) input_mask_gated[127];
  assign vec_sum_002 = vec_sum_001 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:980" *) input_mask_gated[2];
  assign _00609_ = vec_data_000 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13186" *) { mask_d1[0], mask_d1[0], mask_d1[0], mask_d1[0], mask_d1[0], mask_d1[0], mask_d1[0], mask_d1[0] };
  assign _00610_ = vec_data_001 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13196" *) { mask_d1[1], mask_d1[1], mask_d1[1], mask_d1[1], mask_d1[1], mask_d1[1], mask_d1[1], mask_d1[1] };
  assign _00611_ = vec_data_002 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13206" *) { mask_d1[2], mask_d1[2], mask_d1[2], mask_d1[2], mask_d1[2], mask_d1[2], mask_d1[2], mask_d1[2] };
  assign _00612_ = vec_data_003 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13216" *) { mask_d1[3], mask_d1[3], mask_d1[3], mask_d1[3], mask_d1[3], mask_d1[3], mask_d1[3], mask_d1[3] };
  assign _00613_ = vec_data_004 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13226" *) { mask_d1[4], mask_d1[4], mask_d1[4], mask_d1[4], mask_d1[4], mask_d1[4], mask_d1[4], mask_d1[4] };
  assign _00614_ = vec_data_005 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13236" *) { mask_d1[5], mask_d1[5], mask_d1[5], mask_d1[5], mask_d1[5], mask_d1[5], mask_d1[5], mask_d1[5] };
  assign _00615_ = vec_data_006 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13246" *) { mask_d1[6], mask_d1[6], mask_d1[6], mask_d1[6], mask_d1[6], mask_d1[6], mask_d1[6], mask_d1[6] };
  assign _00616_ = vec_data_007 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13256" *) { mask_d1[7], mask_d1[7], mask_d1[7], mask_d1[7], mask_d1[7], mask_d1[7], mask_d1[7], mask_d1[7] };
  assign _00617_ = vec_data_008 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13266" *) { mask_d1[8], mask_d1[8], mask_d1[8], mask_d1[8], mask_d1[8], mask_d1[8], mask_d1[8], mask_d1[8] };
  assign _00618_ = vec_data_009 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13276" *) { mask_d1[9], mask_d1[9], mask_d1[9], mask_d1[9], mask_d1[9], mask_d1[9], mask_d1[9], mask_d1[9] };
  assign _00619_ = vec_data_010 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13286" *) { mask_d1[10], mask_d1[10], mask_d1[10], mask_d1[10], mask_d1[10], mask_d1[10], mask_d1[10], mask_d1[10] };
  assign _00620_ = vec_data_011 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13296" *) { mask_d1[11], mask_d1[11], mask_d1[11], mask_d1[11], mask_d1[11], mask_d1[11], mask_d1[11], mask_d1[11] };
  assign _00621_ = vec_data_012 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13306" *) { mask_d1[12], mask_d1[12], mask_d1[12], mask_d1[12], mask_d1[12], mask_d1[12], mask_d1[12], mask_d1[12] };
  assign _00622_ = vec_data_013 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13316" *) { mask_d1[13], mask_d1[13], mask_d1[13], mask_d1[13], mask_d1[13], mask_d1[13], mask_d1[13], mask_d1[13] };
  assign _00623_ = vec_data_014 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13326" *) { mask_d1[14], mask_d1[14], mask_d1[14], mask_d1[14], mask_d1[14], mask_d1[14], mask_d1[14], mask_d1[14] };
  assign _00624_ = vec_data_015 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13336" *) { mask_d1[15], mask_d1[15], mask_d1[15], mask_d1[15], mask_d1[15], mask_d1[15], mask_d1[15], mask_d1[15] };
  assign _00625_ = vec_data_016 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13346" *) { mask_d1[16], mask_d1[16], mask_d1[16], mask_d1[16], mask_d1[16], mask_d1[16], mask_d1[16], mask_d1[16] };
  assign _00626_ = vec_data_017 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13356" *) { mask_d1[17], mask_d1[17], mask_d1[17], mask_d1[17], mask_d1[17], mask_d1[17], mask_d1[17], mask_d1[17] };
  assign _00627_ = vec_data_018 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13366" *) { mask_d1[18], mask_d1[18], mask_d1[18], mask_d1[18], mask_d1[18], mask_d1[18], mask_d1[18], mask_d1[18] };
  assign _00628_ = vec_data_019 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13376" *) { mask_d1[19], mask_d1[19], mask_d1[19], mask_d1[19], mask_d1[19], mask_d1[19], mask_d1[19], mask_d1[19] };
  assign _00629_ = vec_data_020 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13386" *) { mask_d1[20], mask_d1[20], mask_d1[20], mask_d1[20], mask_d1[20], mask_d1[20], mask_d1[20], mask_d1[20] };
  assign _00630_ = vec_data_021 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13396" *) { mask_d1[21], mask_d1[21], mask_d1[21], mask_d1[21], mask_d1[21], mask_d1[21], mask_d1[21], mask_d1[21] };
  assign _00631_ = vec_data_022 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13406" *) { mask_d1[22], mask_d1[22], mask_d1[22], mask_d1[22], mask_d1[22], mask_d1[22], mask_d1[22], mask_d1[22] };
  assign _00632_ = vec_data_023 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13416" *) { mask_d1[23], mask_d1[23], mask_d1[23], mask_d1[23], mask_d1[23], mask_d1[23], mask_d1[23], mask_d1[23] };
  assign _00633_ = vec_data_024 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13426" *) { mask_d1[24], mask_d1[24], mask_d1[24], mask_d1[24], mask_d1[24], mask_d1[24], mask_d1[24], mask_d1[24] };
  assign _00634_ = vec_data_025 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13436" *) { mask_d1[25], mask_d1[25], mask_d1[25], mask_d1[25], mask_d1[25], mask_d1[25], mask_d1[25], mask_d1[25] };
  assign _00635_ = vec_data_026 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13446" *) { mask_d1[26], mask_d1[26], mask_d1[26], mask_d1[26], mask_d1[26], mask_d1[26], mask_d1[26], mask_d1[26] };
  assign _00636_ = vec_data_027 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13456" *) { mask_d1[27], mask_d1[27], mask_d1[27], mask_d1[27], mask_d1[27], mask_d1[27], mask_d1[27], mask_d1[27] };
  assign _00637_ = vec_data_028 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13466" *) { mask_d1[28], mask_d1[28], mask_d1[28], mask_d1[28], mask_d1[28], mask_d1[28], mask_d1[28], mask_d1[28] };
  assign _00638_ = vec_data_029 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13476" *) { mask_d1[29], mask_d1[29], mask_d1[29], mask_d1[29], mask_d1[29], mask_d1[29], mask_d1[29], mask_d1[29] };
  assign _00639_ = vec_data_030 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13486" *) { mask_d1[30], mask_d1[30], mask_d1[30], mask_d1[30], mask_d1[30], mask_d1[30], mask_d1[30], mask_d1[30] };
  assign _00640_ = vec_data_031 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13496" *) { mask_d1[31], mask_d1[31], mask_d1[31], mask_d1[31], mask_d1[31], mask_d1[31], mask_d1[31], mask_d1[31] };
  assign _00641_ = vec_data_032 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13506" *) { mask_d1[32], mask_d1[32], mask_d1[32], mask_d1[32], mask_d1[32], mask_d1[32], mask_d1[32], mask_d1[32] };
  assign _00642_ = vec_data_033 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13516" *) { mask_d1[33], mask_d1[33], mask_d1[33], mask_d1[33], mask_d1[33], mask_d1[33], mask_d1[33], mask_d1[33] };
  assign _00643_ = vec_data_034 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13526" *) { mask_d1[34], mask_d1[34], mask_d1[34], mask_d1[34], mask_d1[34], mask_d1[34], mask_d1[34], mask_d1[34] };
  assign _00644_ = vec_data_035 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13536" *) { mask_d1[35], mask_d1[35], mask_d1[35], mask_d1[35], mask_d1[35], mask_d1[35], mask_d1[35], mask_d1[35] };
  assign _00645_ = vec_data_036 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13546" *) { mask_d1[36], mask_d1[36], mask_d1[36], mask_d1[36], mask_d1[36], mask_d1[36], mask_d1[36], mask_d1[36] };
  assign _00646_ = vec_data_037 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13556" *) { mask_d1[37], mask_d1[37], mask_d1[37], mask_d1[37], mask_d1[37], mask_d1[37], mask_d1[37], mask_d1[37] };
  assign _00647_ = vec_data_038 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13566" *) { mask_d1[38], mask_d1[38], mask_d1[38], mask_d1[38], mask_d1[38], mask_d1[38], mask_d1[38], mask_d1[38] };
  assign _00648_ = vec_data_039 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13576" *) { mask_d1[39], mask_d1[39], mask_d1[39], mask_d1[39], mask_d1[39], mask_d1[39], mask_d1[39], mask_d1[39] };
  assign _00649_ = vec_data_040 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13586" *) { mask_d1[40], mask_d1[40], mask_d1[40], mask_d1[40], mask_d1[40], mask_d1[40], mask_d1[40], mask_d1[40] };
  assign _00650_ = vec_data_041 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13596" *) { mask_d1[41], mask_d1[41], mask_d1[41], mask_d1[41], mask_d1[41], mask_d1[41], mask_d1[41], mask_d1[41] };
  assign _00651_ = vec_data_042 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13606" *) { mask_d1[42], mask_d1[42], mask_d1[42], mask_d1[42], mask_d1[42], mask_d1[42], mask_d1[42], mask_d1[42] };
  assign _00652_ = vec_data_043 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13616" *) { mask_d1[43], mask_d1[43], mask_d1[43], mask_d1[43], mask_d1[43], mask_d1[43], mask_d1[43], mask_d1[43] };
  assign _00653_ = vec_data_044 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13626" *) { mask_d1[44], mask_d1[44], mask_d1[44], mask_d1[44], mask_d1[44], mask_d1[44], mask_d1[44], mask_d1[44] };
  assign _00654_ = vec_data_045 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13636" *) { mask_d1[45], mask_d1[45], mask_d1[45], mask_d1[45], mask_d1[45], mask_d1[45], mask_d1[45], mask_d1[45] };
  assign _00655_ = vec_data_046 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13646" *) { mask_d1[46], mask_d1[46], mask_d1[46], mask_d1[46], mask_d1[46], mask_d1[46], mask_d1[46], mask_d1[46] };
  assign _00656_ = vec_data_047 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13656" *) { mask_d1[47], mask_d1[47], mask_d1[47], mask_d1[47], mask_d1[47], mask_d1[47], mask_d1[47], mask_d1[47] };
  assign _00657_ = vec_data_048 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13666" *) { mask_d1[48], mask_d1[48], mask_d1[48], mask_d1[48], mask_d1[48], mask_d1[48], mask_d1[48], mask_d1[48] };
  assign _00658_ = vec_data_049 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13676" *) { mask_d1[49], mask_d1[49], mask_d1[49], mask_d1[49], mask_d1[49], mask_d1[49], mask_d1[49], mask_d1[49] };
  assign _00659_ = vec_data_050 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13686" *) { mask_d1[50], mask_d1[50], mask_d1[50], mask_d1[50], mask_d1[50], mask_d1[50], mask_d1[50], mask_d1[50] };
  assign _00660_ = vec_data_051 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13696" *) { mask_d1[51], mask_d1[51], mask_d1[51], mask_d1[51], mask_d1[51], mask_d1[51], mask_d1[51], mask_d1[51] };
  assign _00661_ = vec_data_052 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13706" *) { mask_d1[52], mask_d1[52], mask_d1[52], mask_d1[52], mask_d1[52], mask_d1[52], mask_d1[52], mask_d1[52] };
  assign _00662_ = vec_data_053 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13716" *) { mask_d1[53], mask_d1[53], mask_d1[53], mask_d1[53], mask_d1[53], mask_d1[53], mask_d1[53], mask_d1[53] };
  assign _00663_ = vec_data_054 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13726" *) { mask_d1[54], mask_d1[54], mask_d1[54], mask_d1[54], mask_d1[54], mask_d1[54], mask_d1[54], mask_d1[54] };
  assign _00664_ = vec_data_055 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13736" *) { mask_d1[55], mask_d1[55], mask_d1[55], mask_d1[55], mask_d1[55], mask_d1[55], mask_d1[55], mask_d1[55] };
  assign _00665_ = vec_data_056 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13746" *) { mask_d1[56], mask_d1[56], mask_d1[56], mask_d1[56], mask_d1[56], mask_d1[56], mask_d1[56], mask_d1[56] };
  assign _00666_ = vec_data_057 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13756" *) { mask_d1[57], mask_d1[57], mask_d1[57], mask_d1[57], mask_d1[57], mask_d1[57], mask_d1[57], mask_d1[57] };
  assign _00667_ = vec_data_058 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13766" *) { mask_d1[58], mask_d1[58], mask_d1[58], mask_d1[58], mask_d1[58], mask_d1[58], mask_d1[58], mask_d1[58] };
  assign _00668_ = vec_data_059 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13776" *) { mask_d1[59], mask_d1[59], mask_d1[59], mask_d1[59], mask_d1[59], mask_d1[59], mask_d1[59], mask_d1[59] };
  assign _00669_ = vec_data_060 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13786" *) { mask_d1[60], mask_d1[60], mask_d1[60], mask_d1[60], mask_d1[60], mask_d1[60], mask_d1[60], mask_d1[60] };
  assign _00670_ = vec_data_061 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13796" *) { mask_d1[61], mask_d1[61], mask_d1[61], mask_d1[61], mask_d1[61], mask_d1[61], mask_d1[61], mask_d1[61] };
  assign _00671_ = vec_data_062 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13806" *) { mask_d1[62], mask_d1[62], mask_d1[62], mask_d1[62], mask_d1[62], mask_d1[62], mask_d1[62], mask_d1[62] };
  assign _00672_ = vec_data_063 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13816" *) { mask_d1[63], mask_d1[63], mask_d1[63], mask_d1[63], mask_d1[63], mask_d1[63], mask_d1[63], mask_d1[63] };
  assign _00673_ = vec_data_064 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13826" *) { mask_d1[64], mask_d1[64], mask_d1[64], mask_d1[64], mask_d1[64], mask_d1[64], mask_d1[64], mask_d1[64] };
  assign _00674_ = vec_data_065 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13836" *) { mask_d1[65], mask_d1[65], mask_d1[65], mask_d1[65], mask_d1[65], mask_d1[65], mask_d1[65], mask_d1[65] };
  assign _00675_ = vec_data_066 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13846" *) { mask_d1[66], mask_d1[66], mask_d1[66], mask_d1[66], mask_d1[66], mask_d1[66], mask_d1[66], mask_d1[66] };
  assign _00676_ = vec_data_067 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13856" *) { mask_d1[67], mask_d1[67], mask_d1[67], mask_d1[67], mask_d1[67], mask_d1[67], mask_d1[67], mask_d1[67] };
  assign _00677_ = vec_data_068 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13866" *) { mask_d1[68], mask_d1[68], mask_d1[68], mask_d1[68], mask_d1[68], mask_d1[68], mask_d1[68], mask_d1[68] };
  assign _00678_ = vec_data_069 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13876" *) { mask_d1[69], mask_d1[69], mask_d1[69], mask_d1[69], mask_d1[69], mask_d1[69], mask_d1[69], mask_d1[69] };
  assign _00679_ = vec_data_070 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13886" *) { mask_d1[70], mask_d1[70], mask_d1[70], mask_d1[70], mask_d1[70], mask_d1[70], mask_d1[70], mask_d1[70] };
  assign _00680_ = vec_data_071 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13896" *) { mask_d1[71], mask_d1[71], mask_d1[71], mask_d1[71], mask_d1[71], mask_d1[71], mask_d1[71], mask_d1[71] };
  assign _00681_ = vec_data_072 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13906" *) { mask_d1[72], mask_d1[72], mask_d1[72], mask_d1[72], mask_d1[72], mask_d1[72], mask_d1[72], mask_d1[72] };
  assign _00682_ = vec_data_073 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13916" *) { mask_d1[73], mask_d1[73], mask_d1[73], mask_d1[73], mask_d1[73], mask_d1[73], mask_d1[73], mask_d1[73] };
  assign _00683_ = vec_data_074 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13926" *) { mask_d1[74], mask_d1[74], mask_d1[74], mask_d1[74], mask_d1[74], mask_d1[74], mask_d1[74], mask_d1[74] };
  assign _00684_ = vec_data_075 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13936" *) { mask_d1[75], mask_d1[75], mask_d1[75], mask_d1[75], mask_d1[75], mask_d1[75], mask_d1[75], mask_d1[75] };
  assign _00685_ = vec_data_076 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13946" *) { mask_d1[76], mask_d1[76], mask_d1[76], mask_d1[76], mask_d1[76], mask_d1[76], mask_d1[76], mask_d1[76] };
  assign _00686_ = vec_data_077 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13956" *) { mask_d1[77], mask_d1[77], mask_d1[77], mask_d1[77], mask_d1[77], mask_d1[77], mask_d1[77], mask_d1[77] };
  assign _00687_ = vec_data_078 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13966" *) { mask_d1[78], mask_d1[78], mask_d1[78], mask_d1[78], mask_d1[78], mask_d1[78], mask_d1[78], mask_d1[78] };
  assign _00688_ = vec_data_079 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13976" *) { mask_d1[79], mask_d1[79], mask_d1[79], mask_d1[79], mask_d1[79], mask_d1[79], mask_d1[79], mask_d1[79] };
  assign _00689_ = vec_data_080 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13986" *) { mask_d1[80], mask_d1[80], mask_d1[80], mask_d1[80], mask_d1[80], mask_d1[80], mask_d1[80], mask_d1[80] };
  assign _00690_ = vec_data_081 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13996" *) { mask_d1[81], mask_d1[81], mask_d1[81], mask_d1[81], mask_d1[81], mask_d1[81], mask_d1[81], mask_d1[81] };
  assign _00691_ = vec_data_082 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14006" *) { mask_d1[82], mask_d1[82], mask_d1[82], mask_d1[82], mask_d1[82], mask_d1[82], mask_d1[82], mask_d1[82] };
  assign _00692_ = vec_data_083 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14016" *) { mask_d1[83], mask_d1[83], mask_d1[83], mask_d1[83], mask_d1[83], mask_d1[83], mask_d1[83], mask_d1[83] };
  assign _00693_ = vec_data_084 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14026" *) { mask_d1[84], mask_d1[84], mask_d1[84], mask_d1[84], mask_d1[84], mask_d1[84], mask_d1[84], mask_d1[84] };
  assign _00694_ = vec_data_085 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14036" *) { mask_d1[85], mask_d1[85], mask_d1[85], mask_d1[85], mask_d1[85], mask_d1[85], mask_d1[85], mask_d1[85] };
  assign _00695_ = vec_data_086 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14046" *) { mask_d1[86], mask_d1[86], mask_d1[86], mask_d1[86], mask_d1[86], mask_d1[86], mask_d1[86], mask_d1[86] };
  assign _00696_ = vec_data_087 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14056" *) { mask_d1[87], mask_d1[87], mask_d1[87], mask_d1[87], mask_d1[87], mask_d1[87], mask_d1[87], mask_d1[87] };
  assign _00697_ = vec_data_088 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14066" *) { mask_d1[88], mask_d1[88], mask_d1[88], mask_d1[88], mask_d1[88], mask_d1[88], mask_d1[88], mask_d1[88] };
  assign _00698_ = vec_data_089 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14076" *) { mask_d1[89], mask_d1[89], mask_d1[89], mask_d1[89], mask_d1[89], mask_d1[89], mask_d1[89], mask_d1[89] };
  assign _00699_ = vec_data_090 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14086" *) { mask_d1[90], mask_d1[90], mask_d1[90], mask_d1[90], mask_d1[90], mask_d1[90], mask_d1[90], mask_d1[90] };
  assign _00700_ = vec_data_091 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14096" *) { mask_d1[91], mask_d1[91], mask_d1[91], mask_d1[91], mask_d1[91], mask_d1[91], mask_d1[91], mask_d1[91] };
  assign _00701_ = vec_data_092 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14106" *) { mask_d1[92], mask_d1[92], mask_d1[92], mask_d1[92], mask_d1[92], mask_d1[92], mask_d1[92], mask_d1[92] };
  assign _00702_ = vec_data_093 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14116" *) { mask_d1[93], mask_d1[93], mask_d1[93], mask_d1[93], mask_d1[93], mask_d1[93], mask_d1[93], mask_d1[93] };
  assign _00703_ = vec_data_094 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14126" *) { mask_d1[94], mask_d1[94], mask_d1[94], mask_d1[94], mask_d1[94], mask_d1[94], mask_d1[94], mask_d1[94] };
  assign _00704_ = vec_data_095 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14136" *) { mask_d1[95], mask_d1[95], mask_d1[95], mask_d1[95], mask_d1[95], mask_d1[95], mask_d1[95], mask_d1[95] };
  assign _00705_ = vec_data_096 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14146" *) { mask_d1[96], mask_d1[96], mask_d1[96], mask_d1[96], mask_d1[96], mask_d1[96], mask_d1[96], mask_d1[96] };
  assign _00706_ = vec_data_097 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14156" *) { mask_d1[97], mask_d1[97], mask_d1[97], mask_d1[97], mask_d1[97], mask_d1[97], mask_d1[97], mask_d1[97] };
  assign _00707_ = vec_data_098 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14166" *) { mask_d1[98], mask_d1[98], mask_d1[98], mask_d1[98], mask_d1[98], mask_d1[98], mask_d1[98], mask_d1[98] };
  assign _00708_ = vec_data_099 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14176" *) { mask_d1[99], mask_d1[99], mask_d1[99], mask_d1[99], mask_d1[99], mask_d1[99], mask_d1[99], mask_d1[99] };
  assign _00709_ = vec_data_100 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14186" *) { mask_d1[100], mask_d1[100], mask_d1[100], mask_d1[100], mask_d1[100], mask_d1[100], mask_d1[100], mask_d1[100] };
  assign _00710_ = vec_data_101 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14196" *) { mask_d1[101], mask_d1[101], mask_d1[101], mask_d1[101], mask_d1[101], mask_d1[101], mask_d1[101], mask_d1[101] };
  assign _00711_ = vec_data_102 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14206" *) { mask_d1[102], mask_d1[102], mask_d1[102], mask_d1[102], mask_d1[102], mask_d1[102], mask_d1[102], mask_d1[102] };
  assign _00712_ = vec_data_103 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14216" *) { mask_d1[103], mask_d1[103], mask_d1[103], mask_d1[103], mask_d1[103], mask_d1[103], mask_d1[103], mask_d1[103] };
  assign _00713_ = vec_data_104 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14226" *) { mask_d1[104], mask_d1[104], mask_d1[104], mask_d1[104], mask_d1[104], mask_d1[104], mask_d1[104], mask_d1[104] };
  assign _00714_ = vec_data_105 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14236" *) { mask_d1[105], mask_d1[105], mask_d1[105], mask_d1[105], mask_d1[105], mask_d1[105], mask_d1[105], mask_d1[105] };
  assign _00715_ = vec_data_106 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14246" *) { mask_d1[106], mask_d1[106], mask_d1[106], mask_d1[106], mask_d1[106], mask_d1[106], mask_d1[106], mask_d1[106] };
  assign _00716_ = vec_data_107 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14256" *) { mask_d1[107], mask_d1[107], mask_d1[107], mask_d1[107], mask_d1[107], mask_d1[107], mask_d1[107], mask_d1[107] };
  assign _00717_ = vec_data_108 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14266" *) { mask_d1[108], mask_d1[108], mask_d1[108], mask_d1[108], mask_d1[108], mask_d1[108], mask_d1[108], mask_d1[108] };
  assign _00718_ = vec_data_109 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14276" *) { mask_d1[109], mask_d1[109], mask_d1[109], mask_d1[109], mask_d1[109], mask_d1[109], mask_d1[109], mask_d1[109] };
  assign _00719_ = vec_data_110 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14286" *) { mask_d1[110], mask_d1[110], mask_d1[110], mask_d1[110], mask_d1[110], mask_d1[110], mask_d1[110], mask_d1[110] };
  assign _00720_ = vec_data_111 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14296" *) { mask_d1[111], mask_d1[111], mask_d1[111], mask_d1[111], mask_d1[111], mask_d1[111], mask_d1[111], mask_d1[111] };
  assign _00721_ = vec_data_112 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14306" *) { mask_d1[112], mask_d1[112], mask_d1[112], mask_d1[112], mask_d1[112], mask_d1[112], mask_d1[112], mask_d1[112] };
  assign _00722_ = vec_data_113 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14316" *) { mask_d1[113], mask_d1[113], mask_d1[113], mask_d1[113], mask_d1[113], mask_d1[113], mask_d1[113], mask_d1[113] };
  assign _00723_ = vec_data_114 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14326" *) { mask_d1[114], mask_d1[114], mask_d1[114], mask_d1[114], mask_d1[114], mask_d1[114], mask_d1[114], mask_d1[114] };
  assign _00724_ = vec_data_115 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14336" *) { mask_d1[115], mask_d1[115], mask_d1[115], mask_d1[115], mask_d1[115], mask_d1[115], mask_d1[115], mask_d1[115] };
  assign _00725_ = vec_data_116 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14346" *) { mask_d1[116], mask_d1[116], mask_d1[116], mask_d1[116], mask_d1[116], mask_d1[116], mask_d1[116], mask_d1[116] };
  assign _00726_ = vec_data_117 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14356" *) { mask_d1[117], mask_d1[117], mask_d1[117], mask_d1[117], mask_d1[117], mask_d1[117], mask_d1[117], mask_d1[117] };
  assign _00727_ = vec_data_118 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14366" *) { mask_d1[118], mask_d1[118], mask_d1[118], mask_d1[118], mask_d1[118], mask_d1[118], mask_d1[118], mask_d1[118] };
  assign _00728_ = vec_data_119 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14376" *) { mask_d1[119], mask_d1[119], mask_d1[119], mask_d1[119], mask_d1[119], mask_d1[119], mask_d1[119], mask_d1[119] };
  assign _00729_ = vec_data_120 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14386" *) { mask_d1[120], mask_d1[120], mask_d1[120], mask_d1[120], mask_d1[120], mask_d1[120], mask_d1[120], mask_d1[120] };
  assign _00730_ = vec_data_121 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14396" *) { mask_d1[121], mask_d1[121], mask_d1[121], mask_d1[121], mask_d1[121], mask_d1[121], mask_d1[121], mask_d1[121] };
  assign _00731_ = vec_data_122 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14406" *) { mask_d1[122], mask_d1[122], mask_d1[122], mask_d1[122], mask_d1[122], mask_d1[122], mask_d1[122], mask_d1[122] };
  assign _00732_ = vec_data_123 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14416" *) { mask_d1[123], mask_d1[123], mask_d1[123], mask_d1[123], mask_d1[123], mask_d1[123], mask_d1[123], mask_d1[123] };
  assign _00733_ = vec_data_124 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14426" *) { mask_d1[124], mask_d1[124], mask_d1[124], mask_d1[124], mask_d1[124], mask_d1[124], mask_d1[124], mask_d1[124] };
  assign _00734_ = vec_data_125 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14436" *) { mask_d1[125], mask_d1[125], mask_d1[125], mask_d1[125], mask_d1[125], mask_d1[125], mask_d1[125], mask_d1[125] };
  assign _00735_ = vec_data_126 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14446" *) { mask_d1[126], mask_d1[126], mask_d1[126], mask_d1[126], mask_d1[126], mask_d1[126], mask_d1[126], mask_d1[126] };
  assign _00736_ = vec_data_127 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14456" *) { mask_d1[127], mask_d1[127], mask_d1[127], mask_d1[127], mask_d1[127], mask_d1[127], mask_d1[127], mask_d1[127] };
  assign _00737_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2606" *) input_mask_en[0];
  assign _00738_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2766" *) input_mask_en[1];
  assign _00739_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2926" *) input_mask_en[2];
  assign _00740_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3086" *) input_mask_en[3];
  assign _00741_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3246" *) input_mask_en[4];
  assign _00742_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3406" *) input_mask_en[5];
  assign _00743_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3566" *) input_mask_en[6];
  assign _00744_ = input_pipe_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3726" *) input_mask_en[7];
  always @(posedge nvdla_core_clk)
      vec_data_127_d3 <= _00261_;
  always @(posedge nvdla_core_clk)
      vec_data_126_d3 <= _00259_;
  always @(posedge nvdla_core_clk)
      vec_data_125_d3 <= _00257_;
  always @(posedge nvdla_core_clk)
      vec_data_124_d3 <= _00255_;
  always @(posedge nvdla_core_clk)
      vec_data_123_d3 <= _00253_;
  always @(posedge nvdla_core_clk)
      vec_data_122_d3 <= _00251_;
  always @(posedge nvdla_core_clk)
      vec_data_121_d3 <= _00249_;
  always @(posedge nvdla_core_clk)
      vec_data_120_d3 <= _00247_;
  always @(posedge nvdla_core_clk)
      vec_data_119_d3 <= _00245_;
  always @(posedge nvdla_core_clk)
      vec_data_118_d3 <= _00243_;
  always @(posedge nvdla_core_clk)
      vec_data_117_d3 <= _00241_;
  always @(posedge nvdla_core_clk)
      vec_data_116_d3 <= _00239_;
  always @(posedge nvdla_core_clk)
      vec_data_115_d3 <= _00237_;
  always @(posedge nvdla_core_clk)
      vec_data_114_d3 <= _00235_;
  always @(posedge nvdla_core_clk)
      vec_data_113_d3 <= _00233_;
  always @(posedge nvdla_core_clk)
      vec_data_112_d3 <= _00231_;
  always @(posedge nvdla_core_clk)
      vec_data_111_d3 <= _00229_;
  always @(posedge nvdla_core_clk)
      vec_data_110_d3 <= _00227_;
  always @(posedge nvdla_core_clk)
      vec_data_109_d3 <= _00225_;
  always @(posedge nvdla_core_clk)
      vec_data_108_d3 <= _00223_;
  always @(posedge nvdla_core_clk)
      vec_data_107_d3 <= _00221_;
  always @(posedge nvdla_core_clk)
      vec_data_106_d3 <= _00219_;
  always @(posedge nvdla_core_clk)
      vec_data_105_d3 <= _00217_;
  always @(posedge nvdla_core_clk)
      vec_data_104_d3 <= _00215_;
  always @(posedge nvdla_core_clk)
      vec_data_103_d3 <= _00213_;
  always @(posedge nvdla_core_clk)
      vec_data_102_d3 <= _00211_;
  always @(posedge nvdla_core_clk)
      vec_data_101_d3 <= _00209_;
  always @(posedge nvdla_core_clk)
      vec_data_100_d3 <= _00207_;
  always @(posedge nvdla_core_clk)
      vec_data_099_d3 <= _00205_;
  always @(posedge nvdla_core_clk)
      vec_data_098_d3 <= _00203_;
  always @(posedge nvdla_core_clk)
      vec_data_097_d3 <= _00201_;
  always @(posedge nvdla_core_clk)
      vec_data_096_d3 <= _00199_;
  always @(posedge nvdla_core_clk)
      vec_data_095_d3 <= _00197_;
  always @(posedge nvdla_core_clk)
      vec_data_094_d3 <= _00195_;
  always @(posedge nvdla_core_clk)
      vec_data_093_d3 <= _00193_;
  always @(posedge nvdla_core_clk)
      vec_data_092_d3 <= _00191_;
  always @(posedge nvdla_core_clk)
      vec_data_091_d3 <= _00189_;
  always @(posedge nvdla_core_clk)
      vec_data_090_d3 <= _00187_;
  always @(posedge nvdla_core_clk)
      vec_data_089_d3 <= _00185_;
  always @(posedge nvdla_core_clk)
      vec_data_088_d3 <= _00183_;
  always @(posedge nvdla_core_clk)
      vec_data_087_d3 <= _00181_;
  always @(posedge nvdla_core_clk)
      vec_data_086_d3 <= _00179_;
  always @(posedge nvdla_core_clk)
      vec_data_085_d3 <= _00177_;
  always @(posedge nvdla_core_clk)
      vec_data_084_d3 <= _00175_;
  always @(posedge nvdla_core_clk)
      vec_data_083_d3 <= _00173_;
  always @(posedge nvdla_core_clk)
      vec_data_082_d3 <= _00171_;
  always @(posedge nvdla_core_clk)
      vec_data_081_d3 <= _00169_;
  always @(posedge nvdla_core_clk)
      vec_data_080_d3 <= _00167_;
  always @(posedge nvdla_core_clk)
      vec_data_079_d3 <= _00165_;
  always @(posedge nvdla_core_clk)
      vec_data_078_d3 <= _00163_;
  always @(posedge nvdla_core_clk)
      vec_data_077_d3 <= _00161_;
  always @(posedge nvdla_core_clk)
      vec_data_076_d3 <= _00159_;
  always @(posedge nvdla_core_clk)
      vec_data_075_d3 <= _00157_;
  always @(posedge nvdla_core_clk)
      vec_data_074_d3 <= _00155_;
  always @(posedge nvdla_core_clk)
      vec_data_073_d3 <= _00153_;
  always @(posedge nvdla_core_clk)
      vec_data_072_d3 <= _00151_;
  always @(posedge nvdla_core_clk)
      vec_data_071_d3 <= _00149_;
  always @(posedge nvdla_core_clk)
      vec_data_070_d3 <= _00147_;
  always @(posedge nvdla_core_clk)
      vec_data_069_d3 <= _00145_;
  always @(posedge nvdla_core_clk)
      vec_data_068_d3 <= _00143_;
  always @(posedge nvdla_core_clk)
      vec_data_067_d3 <= _00141_;
  always @(posedge nvdla_core_clk)
      vec_data_066_d3 <= _00139_;
  always @(posedge nvdla_core_clk)
      vec_data_065_d3 <= _00137_;
  always @(posedge nvdla_core_clk)
      vec_data_064_d3 <= _00135_;
  always @(posedge nvdla_core_clk)
      vec_data_063_d3 <= _00133_;
  always @(posedge nvdla_core_clk)
      vec_data_062_d3 <= _00131_;
  always @(posedge nvdla_core_clk)
      vec_data_061_d3 <= _00129_;
  always @(posedge nvdla_core_clk)
      vec_data_060_d3 <= _00127_;
  always @(posedge nvdla_core_clk)
      vec_data_059_d3 <= _00125_;
  always @(posedge nvdla_core_clk)
      vec_data_058_d3 <= _00123_;
  always @(posedge nvdla_core_clk)
      vec_data_057_d3 <= _00121_;
  always @(posedge nvdla_core_clk)
      vec_data_056_d3 <= _00119_;
  always @(posedge nvdla_core_clk)
      vec_data_055_d3 <= _00117_;
  always @(posedge nvdla_core_clk)
      vec_data_054_d3 <= _00115_;
  always @(posedge nvdla_core_clk)
      vec_data_053_d3 <= _00113_;
  always @(posedge nvdla_core_clk)
      vec_data_052_d3 <= _00111_;
  always @(posedge nvdla_core_clk)
      vec_data_051_d3 <= _00109_;
  always @(posedge nvdla_core_clk)
      vec_data_050_d3 <= _00107_;
  always @(posedge nvdla_core_clk)
      vec_data_049_d3 <= _00105_;
  always @(posedge nvdla_core_clk)
      vec_data_048_d3 <= _00103_;
  always @(posedge nvdla_core_clk)
      vec_data_047_d3 <= _00101_;
  always @(posedge nvdla_core_clk)
      vec_data_046_d3 <= _00099_;
  always @(posedge nvdla_core_clk)
      vec_data_045_d3 <= _00097_;
  always @(posedge nvdla_core_clk)
      vec_data_044_d3 <= _00095_;
  always @(posedge nvdla_core_clk)
      vec_data_043_d3 <= _00093_;
  always @(posedge nvdla_core_clk)
      vec_data_042_d3 <= _00091_;
  always @(posedge nvdla_core_clk)
      vec_data_041_d3 <= _00089_;
  always @(posedge nvdla_core_clk)
      vec_data_040_d3 <= _00087_;
  always @(posedge nvdla_core_clk)
      vec_data_039_d3 <= _00085_;
  always @(posedge nvdla_core_clk)
      vec_data_038_d3 <= _00083_;
  always @(posedge nvdla_core_clk)
      vec_data_037_d3 <= _00081_;
  always @(posedge nvdla_core_clk)
      vec_data_036_d3 <= _00079_;
  always @(posedge nvdla_core_clk)
      vec_data_035_d3 <= _00077_;
  always @(posedge nvdla_core_clk)
      vec_data_034_d3 <= _00075_;
  always @(posedge nvdla_core_clk)
      vec_data_033_d3 <= _00073_;
  always @(posedge nvdla_core_clk)
      vec_data_032_d3 <= _00071_;
  always @(posedge nvdla_core_clk)
      vec_data_031_d3 <= _00069_;
  always @(posedge nvdla_core_clk)
      vec_data_030_d3 <= _00067_;
  always @(posedge nvdla_core_clk)
      vec_data_029_d3 <= _00065_;
  always @(posedge nvdla_core_clk)
      vec_data_028_d3 <= _00063_;
  always @(posedge nvdla_core_clk)
      vec_data_027_d3 <= _00061_;
  always @(posedge nvdla_core_clk)
      vec_data_026_d3 <= _00059_;
  always @(posedge nvdla_core_clk)
      vec_data_025_d3 <= _00057_;
  always @(posedge nvdla_core_clk)
      vec_data_024_d3 <= _00055_;
  always @(posedge nvdla_core_clk)
      vec_data_023_d3 <= _00053_;
  always @(posedge nvdla_core_clk)
      vec_data_022_d3 <= _00051_;
  always @(posedge nvdla_core_clk)
      vec_data_021_d3 <= _00049_;
  always @(posedge nvdla_core_clk)
      vec_data_020_d3 <= _00047_;
  always @(posedge nvdla_core_clk)
      vec_data_019_d3 <= _00045_;
  always @(posedge nvdla_core_clk)
      vec_data_018_d3 <= _00043_;
  always @(posedge nvdla_core_clk)
      vec_data_017_d3 <= _00041_;
  always @(posedge nvdla_core_clk)
      vec_data_016_d3 <= _00039_;
  always @(posedge nvdla_core_clk)
      vec_data_015_d3 <= _00037_;
  always @(posedge nvdla_core_clk)
      vec_data_014_d3 <= _00035_;
  always @(posedge nvdla_core_clk)
      vec_data_013_d3 <= _00033_;
  always @(posedge nvdla_core_clk)
      vec_data_012_d3 <= _00031_;
  always @(posedge nvdla_core_clk)
      vec_data_011_d3 <= _00029_;
  always @(posedge nvdla_core_clk)
      vec_data_010_d3 <= _00027_;
  always @(posedge nvdla_core_clk)
      vec_data_009_d3 <= _00025_;
  always @(posedge nvdla_core_clk)
      vec_data_008_d3 <= _00023_;
  always @(posedge nvdla_core_clk)
      vec_data_007_d3 <= _00021_;
  always @(posedge nvdla_core_clk)
      vec_data_006_d3 <= _00019_;
  always @(posedge nvdla_core_clk)
      vec_data_005_d3 <= _00017_;
  always @(posedge nvdla_core_clk)
      vec_data_004_d3 <= _00015_;
  always @(posedge nvdla_core_clk)
      vec_data_003_d3 <= _00013_;
  always @(posedge nvdla_core_clk)
      vec_data_002_d3 <= _00011_;
  always @(posedge nvdla_core_clk)
      vec_data_001_d3 <= _00009_;
  always @(posedge nvdla_core_clk)
      vec_data_000_d3 <= _00007_;
  always @(posedge nvdla_core_clk)
      sel_d3 <= _00005_;
  always @(posedge nvdla_core_clk)
      mask_d3 <= _00002_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      valid_d3 <= 1'b0;
    else
      valid_d3 <= valid_d2;
  always @(posedge nvdla_core_clk)
      vec_data_127_d2 <= _00260_;
  always @(posedge nvdla_core_clk)
      vec_data_126_d2 <= _00258_;
  always @(posedge nvdla_core_clk)
      vec_data_125_d2 <= _00256_;
  always @(posedge nvdla_core_clk)
      vec_data_124_d2 <= _00254_;
  always @(posedge nvdla_core_clk)
      vec_data_123_d2 <= _00252_;
  always @(posedge nvdla_core_clk)
      vec_data_122_d2 <= _00250_;
  always @(posedge nvdla_core_clk)
      vec_data_121_d2 <= _00248_;
  always @(posedge nvdla_core_clk)
      vec_data_120_d2 <= _00246_;
  always @(posedge nvdla_core_clk)
      vec_data_119_d2 <= _00244_;
  always @(posedge nvdla_core_clk)
      vec_data_118_d2 <= _00242_;
  always @(posedge nvdla_core_clk)
      vec_data_117_d2 <= _00240_;
  always @(posedge nvdla_core_clk)
      vec_data_116_d2 <= _00238_;
  always @(posedge nvdla_core_clk)
      vec_data_115_d2 <= _00236_;
  always @(posedge nvdla_core_clk)
      vec_data_114_d2 <= _00234_;
  always @(posedge nvdla_core_clk)
      vec_data_113_d2 <= _00232_;
  always @(posedge nvdla_core_clk)
      vec_data_112_d2 <= _00230_;
  always @(posedge nvdla_core_clk)
      vec_data_111_d2 <= _00228_;
  always @(posedge nvdla_core_clk)
      vec_data_110_d2 <= _00226_;
  always @(posedge nvdla_core_clk)
      vec_data_109_d2 <= _00224_;
  always @(posedge nvdla_core_clk)
      vec_data_108_d2 <= _00222_;
  always @(posedge nvdla_core_clk)
      vec_data_107_d2 <= _00220_;
  always @(posedge nvdla_core_clk)
      vec_data_106_d2 <= _00218_;
  always @(posedge nvdla_core_clk)
      vec_data_105_d2 <= _00216_;
  always @(posedge nvdla_core_clk)
      vec_data_104_d2 <= _00214_;
  always @(posedge nvdla_core_clk)
      vec_data_103_d2 <= _00212_;
  always @(posedge nvdla_core_clk)
      vec_data_102_d2 <= _00210_;
  always @(posedge nvdla_core_clk)
      vec_data_101_d2 <= _00208_;
  always @(posedge nvdla_core_clk)
      vec_data_100_d2 <= _00206_;
  always @(posedge nvdla_core_clk)
      vec_data_099_d2 <= _00204_;
  always @(posedge nvdla_core_clk)
      vec_data_098_d2 <= _00202_;
  always @(posedge nvdla_core_clk)
      vec_data_097_d2 <= _00200_;
  always @(posedge nvdla_core_clk)
      vec_data_096_d2 <= _00198_;
  always @(posedge nvdla_core_clk)
      vec_data_095_d2 <= _00196_;
  always @(posedge nvdla_core_clk)
      vec_data_094_d2 <= _00194_;
  always @(posedge nvdla_core_clk)
      vec_data_093_d2 <= _00192_;
  always @(posedge nvdla_core_clk)
      vec_data_092_d2 <= _00190_;
  always @(posedge nvdla_core_clk)
      vec_data_091_d2 <= _00188_;
  always @(posedge nvdla_core_clk)
      vec_data_090_d2 <= _00186_;
  always @(posedge nvdla_core_clk)
      vec_data_089_d2 <= _00184_;
  always @(posedge nvdla_core_clk)
      vec_data_088_d2 <= _00182_;
  always @(posedge nvdla_core_clk)
      vec_data_087_d2 <= _00180_;
  always @(posedge nvdla_core_clk)
      vec_data_086_d2 <= _00178_;
  always @(posedge nvdla_core_clk)
      vec_data_085_d2 <= _00176_;
  always @(posedge nvdla_core_clk)
      vec_data_084_d2 <= _00174_;
  always @(posedge nvdla_core_clk)
      vec_data_083_d2 <= _00172_;
  always @(posedge nvdla_core_clk)
      vec_data_082_d2 <= _00170_;
  always @(posedge nvdla_core_clk)
      vec_data_081_d2 <= _00168_;
  always @(posedge nvdla_core_clk)
      vec_data_080_d2 <= _00166_;
  always @(posedge nvdla_core_clk)
      vec_data_079_d2 <= _00164_;
  always @(posedge nvdla_core_clk)
      vec_data_078_d2 <= _00162_;
  always @(posedge nvdla_core_clk)
      vec_data_077_d2 <= _00160_;
  always @(posedge nvdla_core_clk)
      vec_data_076_d2 <= _00158_;
  always @(posedge nvdla_core_clk)
      vec_data_075_d2 <= _00156_;
  always @(posedge nvdla_core_clk)
      vec_data_074_d2 <= _00154_;
  always @(posedge nvdla_core_clk)
      vec_data_073_d2 <= _00152_;
  always @(posedge nvdla_core_clk)
      vec_data_072_d2 <= _00150_;
  always @(posedge nvdla_core_clk)
      vec_data_071_d2 <= _00148_;
  always @(posedge nvdla_core_clk)
      vec_data_070_d2 <= _00146_;
  always @(posedge nvdla_core_clk)
      vec_data_069_d2 <= _00144_;
  always @(posedge nvdla_core_clk)
      vec_data_068_d2 <= _00142_;
  always @(posedge nvdla_core_clk)
      vec_data_067_d2 <= _00140_;
  always @(posedge nvdla_core_clk)
      vec_data_066_d2 <= _00138_;
  always @(posedge nvdla_core_clk)
      vec_data_065_d2 <= _00136_;
  always @(posedge nvdla_core_clk)
      vec_data_064_d2 <= _00134_;
  always @(posedge nvdla_core_clk)
      vec_data_063_d2 <= _00132_;
  always @(posedge nvdla_core_clk)
      vec_data_062_d2 <= _00130_;
  always @(posedge nvdla_core_clk)
      vec_data_061_d2 <= _00128_;
  always @(posedge nvdla_core_clk)
      vec_data_060_d2 <= _00126_;
  always @(posedge nvdla_core_clk)
      vec_data_059_d2 <= _00124_;
  always @(posedge nvdla_core_clk)
      vec_data_058_d2 <= _00122_;
  always @(posedge nvdla_core_clk)
      vec_data_057_d2 <= _00120_;
  always @(posedge nvdla_core_clk)
      vec_data_056_d2 <= _00118_;
  always @(posedge nvdla_core_clk)
      vec_data_055_d2 <= _00116_;
  always @(posedge nvdla_core_clk)
      vec_data_054_d2 <= _00114_;
  always @(posedge nvdla_core_clk)
      vec_data_053_d2 <= _00112_;
  always @(posedge nvdla_core_clk)
      vec_data_052_d2 <= _00110_;
  always @(posedge nvdla_core_clk)
      vec_data_051_d2 <= _00108_;
  always @(posedge nvdla_core_clk)
      vec_data_050_d2 <= _00106_;
  always @(posedge nvdla_core_clk)
      vec_data_049_d2 <= _00104_;
  always @(posedge nvdla_core_clk)
      vec_data_048_d2 <= _00102_;
  always @(posedge nvdla_core_clk)
      vec_data_047_d2 <= _00100_;
  always @(posedge nvdla_core_clk)
      vec_data_046_d2 <= _00098_;
  always @(posedge nvdla_core_clk)
      vec_data_045_d2 <= _00096_;
  always @(posedge nvdla_core_clk)
      vec_data_044_d2 <= _00094_;
  always @(posedge nvdla_core_clk)
      vec_data_043_d2 <= _00092_;
  always @(posedge nvdla_core_clk)
      vec_data_042_d2 <= _00090_;
  always @(posedge nvdla_core_clk)
      vec_data_041_d2 <= _00088_;
  always @(posedge nvdla_core_clk)
      vec_data_040_d2 <= _00086_;
  always @(posedge nvdla_core_clk)
      vec_data_039_d2 <= _00084_;
  always @(posedge nvdla_core_clk)
      vec_data_038_d2 <= _00082_;
  always @(posedge nvdla_core_clk)
      vec_data_037_d2 <= _00080_;
  always @(posedge nvdla_core_clk)
      vec_data_036_d2 <= _00078_;
  always @(posedge nvdla_core_clk)
      vec_data_035_d2 <= _00076_;
  always @(posedge nvdla_core_clk)
      vec_data_034_d2 <= _00074_;
  always @(posedge nvdla_core_clk)
      vec_data_033_d2 <= _00072_;
  always @(posedge nvdla_core_clk)
      vec_data_032_d2 <= _00070_;
  always @(posedge nvdla_core_clk)
      vec_data_031_d2 <= _00068_;
  always @(posedge nvdla_core_clk)
      vec_data_030_d2 <= _00066_;
  always @(posedge nvdla_core_clk)
      vec_data_029_d2 <= _00064_;
  always @(posedge nvdla_core_clk)
      vec_data_028_d2 <= _00062_;
  always @(posedge nvdla_core_clk)
      vec_data_027_d2 <= _00060_;
  always @(posedge nvdla_core_clk)
      vec_data_026_d2 <= _00058_;
  always @(posedge nvdla_core_clk)
      vec_data_025_d2 <= _00056_;
  always @(posedge nvdla_core_clk)
      vec_data_024_d2 <= _00054_;
  always @(posedge nvdla_core_clk)
      vec_data_023_d2 <= _00052_;
  always @(posedge nvdla_core_clk)
      vec_data_022_d2 <= _00050_;
  always @(posedge nvdla_core_clk)
      vec_data_021_d2 <= _00048_;
  always @(posedge nvdla_core_clk)
      vec_data_020_d2 <= _00046_;
  always @(posedge nvdla_core_clk)
      vec_data_019_d2 <= _00044_;
  always @(posedge nvdla_core_clk)
      vec_data_018_d2 <= _00042_;
  always @(posedge nvdla_core_clk)
      vec_data_017_d2 <= _00040_;
  always @(posedge nvdla_core_clk)
      vec_data_016_d2 <= _00038_;
  always @(posedge nvdla_core_clk)
      vec_data_015_d2 <= _00036_;
  always @(posedge nvdla_core_clk)
      vec_data_014_d2 <= _00034_;
  always @(posedge nvdla_core_clk)
      vec_data_013_d2 <= _00032_;
  always @(posedge nvdla_core_clk)
      vec_data_012_d2 <= _00030_;
  always @(posedge nvdla_core_clk)
      vec_data_011_d2 <= _00028_;
  always @(posedge nvdla_core_clk)
      vec_data_010_d2 <= _00026_;
  always @(posedge nvdla_core_clk)
      vec_data_009_d2 <= _00024_;
  always @(posedge nvdla_core_clk)
      vec_data_008_d2 <= _00022_;
  always @(posedge nvdla_core_clk)
      vec_data_007_d2 <= _00020_;
  always @(posedge nvdla_core_clk)
      vec_data_006_d2 <= _00018_;
  always @(posedge nvdla_core_clk)
      vec_data_005_d2 <= _00016_;
  always @(posedge nvdla_core_clk)
      vec_data_004_d2 <= _00014_;
  always @(posedge nvdla_core_clk)
      vec_data_003_d2 <= _00012_;
  always @(posedge nvdla_core_clk)
      vec_data_002_d2 <= _00010_;
  always @(posedge nvdla_core_clk)
      vec_data_001_d2 <= _00008_;
  always @(posedge nvdla_core_clk)
      vec_data_000_d2 <= _00006_;
  always @(posedge nvdla_core_clk)
      sel_d2 <= _00004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      valid_d2 <= 1'b0;
    else
      valid_d2 <= valid_d1;
  reg [7:0] _09745_;
  always @(posedge nvdla_core_clk)
      _09745_ <= _00389_;
  assign { _00745_[7], vec_sum_127_d1 } = _09745_;
  always @(posedge nvdla_core_clk)
      vec_sum_126_d1 <= _00388_;
  always @(posedge nvdla_core_clk)
      vec_sum_125_d1 <= _00387_;
  always @(posedge nvdla_core_clk)
      vec_sum_124_d1 <= _00386_;
  always @(posedge nvdla_core_clk)
      vec_sum_123_d1 <= _00385_;
  always @(posedge nvdla_core_clk)
      vec_sum_122_d1 <= _00384_;
  always @(posedge nvdla_core_clk)
      vec_sum_121_d1 <= _00383_;
  always @(posedge nvdla_core_clk)
      vec_sum_120_d1 <= _00382_;
  always @(posedge nvdla_core_clk)
      vec_sum_119_d1 <= _00381_;
  always @(posedge nvdla_core_clk)
      vec_sum_118_d1 <= _00380_;
  always @(posedge nvdla_core_clk)
      vec_sum_117_d1 <= _00379_;
  always @(posedge nvdla_core_clk)
      vec_sum_116_d1 <= _00378_;
  always @(posedge nvdla_core_clk)
      vec_sum_115_d1 <= _00377_;
  always @(posedge nvdla_core_clk)
      vec_sum_114_d1 <= _00376_;
  always @(posedge nvdla_core_clk)
      vec_sum_113_d1 <= _00375_;
  always @(posedge nvdla_core_clk)
      vec_sum_112_d1 <= _00374_;
  always @(posedge nvdla_core_clk)
      vec_sum_111_d1 <= _00373_;
  always @(posedge nvdla_core_clk)
      vec_sum_110_d1 <= _00372_;
  always @(posedge nvdla_core_clk)
      vec_sum_109_d1 <= _00371_;
  always @(posedge nvdla_core_clk)
      vec_sum_108_d1 <= _00370_;
  always @(posedge nvdla_core_clk)
      vec_sum_107_d1 <= _00369_;
  always @(posedge nvdla_core_clk)
      vec_sum_106_d1 <= _00368_;
  always @(posedge nvdla_core_clk)
      vec_sum_105_d1 <= _00367_;
  always @(posedge nvdla_core_clk)
      vec_sum_104_d1 <= _00366_;
  always @(posedge nvdla_core_clk)
      vec_sum_103_d1 <= _00365_;
  always @(posedge nvdla_core_clk)
      vec_sum_102_d1 <= _00364_;
  always @(posedge nvdla_core_clk)
      vec_sum_101_d1 <= _00363_;
  always @(posedge nvdla_core_clk)
      vec_sum_100_d1 <= _00362_;
  always @(posedge nvdla_core_clk)
      vec_sum_099_d1 <= _00361_;
  always @(posedge nvdla_core_clk)
      vec_sum_098_d1 <= _00360_;
  always @(posedge nvdla_core_clk)
      vec_sum_097_d1 <= _00359_;
  always @(posedge nvdla_core_clk)
      vec_sum_096_d1 <= _00358_;
  always @(posedge nvdla_core_clk)
      vec_sum_095_d1 <= _00357_;
  always @(posedge nvdla_core_clk)
      vec_sum_094_d1 <= _00356_;
  always @(posedge nvdla_core_clk)
      vec_sum_093_d1 <= _00355_;
  always @(posedge nvdla_core_clk)
      vec_sum_092_d1 <= _00354_;
  always @(posedge nvdla_core_clk)
      vec_sum_091_d1 <= _00353_;
  always @(posedge nvdla_core_clk)
      vec_sum_090_d1 <= _00352_;
  always @(posedge nvdla_core_clk)
      vec_sum_089_d1 <= _00351_;
  always @(posedge nvdla_core_clk)
      vec_sum_088_d1 <= _00350_;
  always @(posedge nvdla_core_clk)
      vec_sum_087_d1 <= _00349_;
  always @(posedge nvdla_core_clk)
      vec_sum_086_d1 <= _00348_;
  always @(posedge nvdla_core_clk)
      vec_sum_085_d1 <= _00347_;
  always @(posedge nvdla_core_clk)
      vec_sum_084_d1 <= _00346_;
  always @(posedge nvdla_core_clk)
      vec_sum_083_d1 <= _00345_;
  always @(posedge nvdla_core_clk)
      vec_sum_082_d1 <= _00344_;
  always @(posedge nvdla_core_clk)
      vec_sum_081_d1 <= _00343_;
  always @(posedge nvdla_core_clk)
      vec_sum_080_d1 <= _00342_;
  always @(posedge nvdla_core_clk)
      vec_sum_079_d1 <= _00341_;
  always @(posedge nvdla_core_clk)
      vec_sum_078_d1 <= _00340_;
  always @(posedge nvdla_core_clk)
      vec_sum_077_d1 <= _00339_;
  always @(posedge nvdla_core_clk)
      vec_sum_076_d1 <= _00338_;
  always @(posedge nvdla_core_clk)
      vec_sum_075_d1 <= _00337_;
  always @(posedge nvdla_core_clk)
      vec_sum_074_d1 <= _00336_;
  always @(posedge nvdla_core_clk)
      vec_sum_073_d1 <= _00335_;
  always @(posedge nvdla_core_clk)
      vec_sum_072_d1 <= _00334_;
  always @(posedge nvdla_core_clk)
      vec_sum_071_d1 <= _00333_;
  always @(posedge nvdla_core_clk)
      vec_sum_070_d1 <= _00332_;
  always @(posedge nvdla_core_clk)
      vec_sum_069_d1 <= _00331_;
  always @(posedge nvdla_core_clk)
      vec_sum_068_d1 <= _00330_;
  always @(posedge nvdla_core_clk)
      vec_sum_067_d1 <= _00329_;
  always @(posedge nvdla_core_clk)
      vec_sum_066_d1 <= _00328_;
  always @(posedge nvdla_core_clk)
      vec_sum_065_d1 <= _00327_;
  always @(posedge nvdla_core_clk)
      vec_sum_064_d1 <= _00326_;
  always @(posedge nvdla_core_clk)
      vec_sum_063_d1 <= _00325_;
  always @(posedge nvdla_core_clk)
      vec_sum_062_d1 <= _00324_;
  always @(posedge nvdla_core_clk)
      vec_sum_061_d1 <= _00323_;
  always @(posedge nvdla_core_clk)
      vec_sum_060_d1 <= _00322_;
  always @(posedge nvdla_core_clk)
      vec_sum_059_d1 <= _00321_;
  always @(posedge nvdla_core_clk)
      vec_sum_058_d1 <= _00320_;
  always @(posedge nvdla_core_clk)
      vec_sum_057_d1 <= _00319_;
  always @(posedge nvdla_core_clk)
      vec_sum_056_d1 <= _00318_;
  always @(posedge nvdla_core_clk)
      vec_sum_055_d1 <= _00317_;
  always @(posedge nvdla_core_clk)
      vec_sum_054_d1 <= _00316_;
  always @(posedge nvdla_core_clk)
      vec_sum_053_d1 <= _00315_;
  always @(posedge nvdla_core_clk)
      vec_sum_052_d1 <= _00314_;
  always @(posedge nvdla_core_clk)
      vec_sum_051_d1 <= _00313_;
  always @(posedge nvdla_core_clk)
      vec_sum_050_d1 <= _00312_;
  always @(posedge nvdla_core_clk)
      vec_sum_049_d1 <= _00311_;
  always @(posedge nvdla_core_clk)
      vec_sum_048_d1 <= _00310_;
  always @(posedge nvdla_core_clk)
      vec_sum_047_d1 <= _00309_;
  always @(posedge nvdla_core_clk)
      vec_sum_046_d1 <= _00308_;
  always @(posedge nvdla_core_clk)
      vec_sum_045_d1 <= _00307_;
  always @(posedge nvdla_core_clk)
      vec_sum_044_d1 <= _00306_;
  always @(posedge nvdla_core_clk)
      vec_sum_043_d1 <= _00305_;
  always @(posedge nvdla_core_clk)
      vec_sum_042_d1 <= _00304_;
  always @(posedge nvdla_core_clk)
      vec_sum_041_d1 <= _00303_;
  always @(posedge nvdla_core_clk)
      vec_sum_040_d1 <= _00302_;
  always @(posedge nvdla_core_clk)
      vec_sum_039_d1 <= _00301_;
  always @(posedge nvdla_core_clk)
      vec_sum_038_d1 <= _00300_;
  always @(posedge nvdla_core_clk)
      vec_sum_037_d1 <= _00299_;
  always @(posedge nvdla_core_clk)
      vec_sum_036_d1 <= _00298_;
  always @(posedge nvdla_core_clk)
      vec_sum_035_d1 <= _00297_;
  always @(posedge nvdla_core_clk)
      vec_sum_034_d1 <= _00296_;
  always @(posedge nvdla_core_clk)
      vec_sum_033_d1 <= _00295_;
  always @(posedge nvdla_core_clk)
      vec_sum_032_d1 <= _00294_;
  always @(posedge nvdla_core_clk)
      vec_sum_031_d1 <= _00293_;
  always @(posedge nvdla_core_clk)
      vec_sum_030_d1 <= _00292_;
  always @(posedge nvdla_core_clk)
      vec_sum_029_d1 <= _00291_;
  always @(posedge nvdla_core_clk)
      vec_sum_028_d1 <= _00290_;
  always @(posedge nvdla_core_clk)
      vec_sum_027_d1 <= _00289_;
  always @(posedge nvdla_core_clk)
      vec_sum_026_d1 <= _00288_;
  always @(posedge nvdla_core_clk)
      vec_sum_025_d1 <= _00287_;
  always @(posedge nvdla_core_clk)
      vec_sum_024_d1 <= _00286_;
  always @(posedge nvdla_core_clk)
      vec_sum_023_d1 <= _00285_;
  always @(posedge nvdla_core_clk)
      vec_sum_022_d1 <= _00284_;
  always @(posedge nvdla_core_clk)
      vec_sum_021_d1 <= _00283_;
  always @(posedge nvdla_core_clk)
      vec_sum_020_d1 <= _00282_;
  always @(posedge nvdla_core_clk)
      vec_sum_019_d1 <= _00281_;
  always @(posedge nvdla_core_clk)
      vec_sum_018_d1 <= _00280_;
  always @(posedge nvdla_core_clk)
      vec_sum_017_d1 <= _00279_;
  always @(posedge nvdla_core_clk)
      vec_sum_016_d1 <= _00278_;
  always @(posedge nvdla_core_clk)
      vec_sum_015_d1 <= _00277_;
  always @(posedge nvdla_core_clk)
      vec_sum_014_d1 <= _00276_;
  always @(posedge nvdla_core_clk)
      vec_sum_013_d1 <= _00275_;
  always @(posedge nvdla_core_clk)
      vec_sum_012_d1 <= _00274_;
  always @(posedge nvdla_core_clk)
      vec_sum_011_d1 <= _00273_;
  always @(posedge nvdla_core_clk)
      vec_sum_010_d1 <= _00272_;
  always @(posedge nvdla_core_clk)
      vec_sum_009_d1 <= _00271_;
  always @(posedge nvdla_core_clk)
      vec_sum_008_d1 <= _00270_;
  always @(posedge nvdla_core_clk)
      vec_sum_007_d1 <= _00269_;
  always @(posedge nvdla_core_clk)
      vec_sum_006_d1 <= _00268_;
  always @(posedge nvdla_core_clk)
      vec_sum_005_d1 <= _00267_;
  always @(posedge nvdla_core_clk)
      vec_sum_004_d1 <= _00266_;
  always @(posedge nvdla_core_clk)
      vec_sum_003_d1 <= _00265_;
  always @(posedge nvdla_core_clk)
      vec_sum_002_d1 <= _00264_;
  always @(posedge nvdla_core_clk)
      vec_sum_001_d1 <= _00263_;
  always @(posedge nvdla_core_clk)
      vec_sum_000_d1 <= _00262_;
  always @(posedge nvdla_core_clk)
      sel_d1 <= _00003_;
  always @(posedge nvdla_core_clk)
      mask_d1 <= _00001_;
  always @(posedge nvdla_core_clk)
      data_d1 <= _00000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      valid_d1 <= 1'b0;
    else
      valid_d1 <= input_pipe_valid;
  assign _00261_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22439" *) vec_data_127_d2 : vec_data_127_d3;
  assign _00259_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22429" *) vec_data_126_d2 : vec_data_126_d3;
  assign _00257_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22419" *) vec_data_125_d2 : vec_data_125_d3;
  assign _00255_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22409" *) vec_data_124_d2 : vec_data_124_d3;
  assign _00253_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22399" *) vec_data_123_d2 : vec_data_123_d3;
  assign _00251_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22389" *) vec_data_122_d2 : vec_data_122_d3;
  assign _00249_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22379" *) vec_data_121_d2 : vec_data_121_d3;
  assign _00247_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22369" *) vec_data_120_d2 : vec_data_120_d3;
  assign _00245_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22359" *) vec_data_119_d2 : vec_data_119_d3;
  assign _00243_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22349" *) vec_data_118_d2 : vec_data_118_d3;
  assign _00241_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22339" *) vec_data_117_d2 : vec_data_117_d3;
  assign _00239_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22329" *) vec_data_116_d2 : vec_data_116_d3;
  assign _00237_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22319" *) vec_data_115_d2 : vec_data_115_d3;
  assign _00235_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22309" *) vec_data_114_d2 : vec_data_114_d3;
  assign _00233_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22299" *) vec_data_113_d2 : vec_data_113_d3;
  assign _00231_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22289" *) vec_data_112_d2 : vec_data_112_d3;
  assign _00229_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22279" *) vec_data_111_d2 : vec_data_111_d3;
  assign _00227_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22269" *) vec_data_110_d2 : vec_data_110_d3;
  assign _00225_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22259" *) vec_data_109_d2 : vec_data_109_d3;
  assign _00223_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22249" *) vec_data_108_d2 : vec_data_108_d3;
  assign _00221_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22239" *) vec_data_107_d2 : vec_data_107_d3;
  assign _00219_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22229" *) vec_data_106_d2 : vec_data_106_d3;
  assign _00217_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22219" *) vec_data_105_d2 : vec_data_105_d3;
  assign _00215_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22209" *) vec_data_104_d2 : vec_data_104_d3;
  assign _00213_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22199" *) vec_data_103_d2 : vec_data_103_d3;
  assign _00211_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22189" *) vec_data_102_d2 : vec_data_102_d3;
  assign _00209_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22179" *) vec_data_101_d2 : vec_data_101_d3;
  assign _00207_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22169" *) vec_data_100_d2 : vec_data_100_d3;
  assign _00205_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22159" *) vec_data_099_d2 : vec_data_099_d3;
  assign _00203_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22149" *) vec_data_098_d2 : vec_data_098_d3;
  assign _00201_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22139" *) vec_data_097_d2 : vec_data_097_d3;
  assign _00199_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22129" *) vec_data_096_d2 : vec_data_096_d3;
  assign _00197_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22119" *) vec_data_095_d2 : vec_data_095_d3;
  assign _00195_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22109" *) vec_data_094_d2 : vec_data_094_d3;
  assign _00193_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22099" *) vec_data_093_d2 : vec_data_093_d3;
  assign _00191_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22089" *) vec_data_092_d2 : vec_data_092_d3;
  assign _00189_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22079" *) vec_data_091_d2 : vec_data_091_d3;
  assign _00187_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22069" *) vec_data_090_d2 : vec_data_090_d3;
  assign _00185_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22059" *) vec_data_089_d2 : vec_data_089_d3;
  assign _00183_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22049" *) vec_data_088_d2 : vec_data_088_d3;
  assign _00181_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22039" *) vec_data_087_d2 : vec_data_087_d3;
  assign _00179_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22029" *) vec_data_086_d2 : vec_data_086_d3;
  assign _00177_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22019" *) vec_data_085_d2 : vec_data_085_d3;
  assign _00175_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:22009" *) vec_data_084_d2 : vec_data_084_d3;
  assign _00173_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21999" *) vec_data_083_d2 : vec_data_083_d3;
  assign _00171_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21989" *) vec_data_082_d2 : vec_data_082_d3;
  assign _00169_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21979" *) vec_data_081_d2 : vec_data_081_d3;
  assign _00167_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21969" *) vec_data_080_d2 : vec_data_080_d3;
  assign _00165_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21959" *) vec_data_079_d2 : vec_data_079_d3;
  assign _00163_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21949" *) vec_data_078_d2 : vec_data_078_d3;
  assign _00161_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21939" *) vec_data_077_d2 : vec_data_077_d3;
  assign _00159_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21929" *) vec_data_076_d2 : vec_data_076_d3;
  assign _00157_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21919" *) vec_data_075_d2 : vec_data_075_d3;
  assign _00155_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21909" *) vec_data_074_d2 : vec_data_074_d3;
  assign _00153_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21899" *) vec_data_073_d2 : vec_data_073_d3;
  assign _00151_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21889" *) vec_data_072_d2 : vec_data_072_d3;
  assign _00149_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21879" *) vec_data_071_d2 : vec_data_071_d3;
  assign _00147_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21869" *) vec_data_070_d2 : vec_data_070_d3;
  assign _00145_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21859" *) vec_data_069_d2 : vec_data_069_d3;
  assign _00143_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21849" *) vec_data_068_d2 : vec_data_068_d3;
  assign _00141_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21839" *) vec_data_067_d2 : vec_data_067_d3;
  assign _00139_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21829" *) vec_data_066_d2 : vec_data_066_d3;
  assign _00137_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21819" *) vec_data_065_d2 : vec_data_065_d3;
  assign _00135_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21809" *) vec_data_064_d2 : vec_data_064_d3;
  assign _00133_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21799" *) vec_data_063_d2 : vec_data_063_d3;
  assign _00131_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21789" *) vec_data_062_d2 : vec_data_062_d3;
  assign _00129_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21779" *) vec_data_061_d2 : vec_data_061_d3;
  assign _00127_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21769" *) vec_data_060_d2 : vec_data_060_d3;
  assign _00125_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21759" *) vec_data_059_d2 : vec_data_059_d3;
  assign _00123_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21749" *) vec_data_058_d2 : vec_data_058_d3;
  assign _00121_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21739" *) vec_data_057_d2 : vec_data_057_d3;
  assign _00119_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21729" *) vec_data_056_d2 : vec_data_056_d3;
  assign _00117_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21719" *) vec_data_055_d2 : vec_data_055_d3;
  assign _00115_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21709" *) vec_data_054_d2 : vec_data_054_d3;
  assign _00113_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21699" *) vec_data_053_d2 : vec_data_053_d3;
  assign _00111_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21689" *) vec_data_052_d2 : vec_data_052_d3;
  assign _00109_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21679" *) vec_data_051_d2 : vec_data_051_d3;
  assign _00107_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21669" *) vec_data_050_d2 : vec_data_050_d3;
  assign _00105_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21659" *) vec_data_049_d2 : vec_data_049_d3;
  assign _00103_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21649" *) vec_data_048_d2 : vec_data_048_d3;
  assign _00101_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21639" *) vec_data_047_d2 : vec_data_047_d3;
  assign _00099_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21629" *) vec_data_046_d2 : vec_data_046_d3;
  assign _00097_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21619" *) vec_data_045_d2 : vec_data_045_d3;
  assign _00095_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21609" *) vec_data_044_d2 : vec_data_044_d3;
  assign _00093_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21599" *) vec_data_043_d2 : vec_data_043_d3;
  assign _00091_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21589" *) vec_data_042_d2 : vec_data_042_d3;
  assign _00089_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21579" *) vec_data_041_d2 : vec_data_041_d3;
  assign _00087_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21569" *) vec_data_040_d2 : vec_data_040_d3;
  assign _00085_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21559" *) vec_data_039_d2 : vec_data_039_d3;
  assign _00083_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21549" *) vec_data_038_d2 : vec_data_038_d3;
  assign _00081_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21539" *) vec_data_037_d2 : vec_data_037_d3;
  assign _00079_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21529" *) vec_data_036_d2 : vec_data_036_d3;
  assign _00077_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21519" *) vec_data_035_d2 : vec_data_035_d3;
  assign _00075_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21509" *) vec_data_034_d2 : vec_data_034_d3;
  assign _00073_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21499" *) vec_data_033_d2 : vec_data_033_d3;
  assign _00071_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21489" *) vec_data_032_d2 : vec_data_032_d3;
  assign _00069_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21479" *) vec_data_031_d2 : vec_data_031_d3;
  assign _00067_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21469" *) vec_data_030_d2 : vec_data_030_d3;
  assign _00065_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21459" *) vec_data_029_d2 : vec_data_029_d3;
  assign _00063_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21449" *) vec_data_028_d2 : vec_data_028_d3;
  assign _00061_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21439" *) vec_data_027_d2 : vec_data_027_d3;
  assign _00059_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21429" *) vec_data_026_d2 : vec_data_026_d3;
  assign _00057_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21419" *) vec_data_025_d2 : vec_data_025_d3;
  assign _00055_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21409" *) vec_data_024_d2 : vec_data_024_d3;
  assign _00053_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21399" *) vec_data_023_d2 : vec_data_023_d3;
  assign _00051_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21389" *) vec_data_022_d2 : vec_data_022_d3;
  assign _00049_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21379" *) vec_data_021_d2 : vec_data_021_d3;
  assign _00047_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21369" *) vec_data_020_d2 : vec_data_020_d3;
  assign _00045_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21359" *) vec_data_019_d2 : vec_data_019_d3;
  assign _00043_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21349" *) vec_data_018_d2 : vec_data_018_d3;
  assign _00041_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21339" *) vec_data_017_d2 : vec_data_017_d3;
  assign _00039_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21329" *) vec_data_016_d2 : vec_data_016_d3;
  assign _00037_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21319" *) vec_data_015_d2 : vec_data_015_d3;
  assign _00035_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21309" *) vec_data_014_d2 : vec_data_014_d3;
  assign _00033_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21299" *) vec_data_013_d2 : vec_data_013_d3;
  assign _00031_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21289" *) vec_data_012_d2 : vec_data_012_d3;
  assign _00029_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21279" *) vec_data_011_d2 : vec_data_011_d3;
  assign _00027_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21269" *) vec_data_010_d2 : vec_data_010_d3;
  assign _00025_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21259" *) vec_data_009_d2 : vec_data_009_d3;
  assign _00023_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21249" *) vec_data_008_d2 : vec_data_008_d3;
  assign _00021_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21239" *) vec_data_007_d2 : vec_data_007_d3;
  assign _00019_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21229" *) vec_data_006_d2 : vec_data_006_d3;
  assign _00017_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21219" *) vec_data_005_d2 : vec_data_005_d3;
  assign _00015_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21209" *) vec_data_004_d2 : vec_data_004_d3;
  assign _00013_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21199" *) vec_data_003_d2 : vec_data_003_d3;
  assign _00011_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21189" *) vec_data_002_d2 : vec_data_002_d3;
  assign _00009_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21179" *) vec_data_001_d2 : vec_data_001_d3;
  assign _00007_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21169" *) vec_data_000_d2 : vec_data_000_d3;
  assign _00005_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21159" *) sel_d2 : sel_d3;
  assign _00002_ = valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21149" *) mask_d2_w : mask_d3;
  assign _00260_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14455" *) _00736_ : vec_data_127_d2;
  assign _00258_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14445" *) _00735_ : vec_data_126_d2;
  assign _00256_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14435" *) _00734_ : vec_data_125_d2;
  assign _00254_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14425" *) _00733_ : vec_data_124_d2;
  assign _00252_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14415" *) _00732_ : vec_data_123_d2;
  assign _00250_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14405" *) _00731_ : vec_data_122_d2;
  assign _00248_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14395" *) _00730_ : vec_data_121_d2;
  assign _00246_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14385" *) _00729_ : vec_data_120_d2;
  assign _00244_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14375" *) _00728_ : vec_data_119_d2;
  assign _00242_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14365" *) _00727_ : vec_data_118_d2;
  assign _00240_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14355" *) _00726_ : vec_data_117_d2;
  assign _00238_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14345" *) _00725_ : vec_data_116_d2;
  assign _00236_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14335" *) _00724_ : vec_data_115_d2;
  assign _00234_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14325" *) _00723_ : vec_data_114_d2;
  assign _00232_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14315" *) _00722_ : vec_data_113_d2;
  assign _00230_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14305" *) _00721_ : vec_data_112_d2;
  assign _00228_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14295" *) _00720_ : vec_data_111_d2;
  assign _00226_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14285" *) _00719_ : vec_data_110_d2;
  assign _00224_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14275" *) _00718_ : vec_data_109_d2;
  assign _00222_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14265" *) _00717_ : vec_data_108_d2;
  assign _00220_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14255" *) _00716_ : vec_data_107_d2;
  assign _00218_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14245" *) _00715_ : vec_data_106_d2;
  assign _00216_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14235" *) _00714_ : vec_data_105_d2;
  assign _00214_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14225" *) _00713_ : vec_data_104_d2;
  assign _00212_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14215" *) _00712_ : vec_data_103_d2;
  assign _00210_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14205" *) _00711_ : vec_data_102_d2;
  assign _00208_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14195" *) _00710_ : vec_data_101_d2;
  assign _00206_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14185" *) _00709_ : vec_data_100_d2;
  assign _00204_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14175" *) _00708_ : vec_data_099_d2;
  assign _00202_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14165" *) _00707_ : vec_data_098_d2;
  assign _00200_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14155" *) _00706_ : vec_data_097_d2;
  assign _00198_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14145" *) _00705_ : vec_data_096_d2;
  assign _00196_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14135" *) _00704_ : vec_data_095_d2;
  assign _00194_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14125" *) _00703_ : vec_data_094_d2;
  assign _00192_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14115" *) _00702_ : vec_data_093_d2;
  assign _00190_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14105" *) _00701_ : vec_data_092_d2;
  assign _00188_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14095" *) _00700_ : vec_data_091_d2;
  assign _00186_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14085" *) _00699_ : vec_data_090_d2;
  assign _00184_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14075" *) _00698_ : vec_data_089_d2;
  assign _00182_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14065" *) _00697_ : vec_data_088_d2;
  assign _00180_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14055" *) _00696_ : vec_data_087_d2;
  assign _00178_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14045" *) _00695_ : vec_data_086_d2;
  assign _00176_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14035" *) _00694_ : vec_data_085_d2;
  assign _00174_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14025" *) _00693_ : vec_data_084_d2;
  assign _00172_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14015" *) _00692_ : vec_data_083_d2;
  assign _00170_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:14005" *) _00691_ : vec_data_082_d2;
  assign _00168_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13995" *) _00690_ : vec_data_081_d2;
  assign _00166_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13985" *) _00689_ : vec_data_080_d2;
  assign _00164_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13975" *) _00688_ : vec_data_079_d2;
  assign _00162_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13965" *) _00687_ : vec_data_078_d2;
  assign _00160_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13955" *) _00686_ : vec_data_077_d2;
  assign _00158_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13945" *) _00685_ : vec_data_076_d2;
  assign _00156_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13935" *) _00684_ : vec_data_075_d2;
  assign _00154_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13925" *) _00683_ : vec_data_074_d2;
  assign _00152_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13915" *) _00682_ : vec_data_073_d2;
  assign _00150_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13905" *) _00681_ : vec_data_072_d2;
  assign _00148_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13895" *) _00680_ : vec_data_071_d2;
  assign _00146_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13885" *) _00679_ : vec_data_070_d2;
  assign _00144_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13875" *) _00678_ : vec_data_069_d2;
  assign _00142_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13865" *) _00677_ : vec_data_068_d2;
  assign _00140_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13855" *) _00676_ : vec_data_067_d2;
  assign _00138_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13845" *) _00675_ : vec_data_066_d2;
  assign _00136_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13835" *) _00674_ : vec_data_065_d2;
  assign _00134_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13825" *) _00673_ : vec_data_064_d2;
  assign _00132_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13815" *) _00672_ : vec_data_063_d2;
  assign _00130_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13805" *) _00671_ : vec_data_062_d2;
  assign _00128_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13795" *) _00670_ : vec_data_061_d2;
  assign _00126_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13785" *) _00669_ : vec_data_060_d2;
  assign _00124_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13775" *) _00668_ : vec_data_059_d2;
  assign _00122_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13765" *) _00667_ : vec_data_058_d2;
  assign _00120_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13755" *) _00666_ : vec_data_057_d2;
  assign _00118_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13745" *) _00665_ : vec_data_056_d2;
  assign _00116_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13735" *) _00664_ : vec_data_055_d2;
  assign _00114_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13725" *) _00663_ : vec_data_054_d2;
  assign _00112_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13715" *) _00662_ : vec_data_053_d2;
  assign _00110_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13705" *) _00661_ : vec_data_052_d2;
  assign _00108_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13695" *) _00660_ : vec_data_051_d2;
  assign _00106_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13685" *) _00659_ : vec_data_050_d2;
  assign _00104_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13675" *) _00658_ : vec_data_049_d2;
  assign _00102_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13665" *) _00657_ : vec_data_048_d2;
  assign _00100_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13655" *) _00656_ : vec_data_047_d2;
  assign _00098_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13645" *) _00655_ : vec_data_046_d2;
  assign _00096_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13635" *) _00654_ : vec_data_045_d2;
  assign _00094_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13625" *) _00653_ : vec_data_044_d2;
  assign _00092_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13615" *) _00652_ : vec_data_043_d2;
  assign _00090_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13605" *) _00651_ : vec_data_042_d2;
  assign _00088_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13595" *) _00650_ : vec_data_041_d2;
  assign _00086_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13585" *) _00649_ : vec_data_040_d2;
  assign _00084_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13575" *) _00648_ : vec_data_039_d2;
  assign _00082_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13565" *) _00647_ : vec_data_038_d2;
  assign _00080_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13555" *) _00646_ : vec_data_037_d2;
  assign _00078_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13545" *) _00645_ : vec_data_036_d2;
  assign _00076_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13535" *) _00644_ : vec_data_035_d2;
  assign _00074_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13525" *) _00643_ : vec_data_034_d2;
  assign _00072_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13515" *) _00642_ : vec_data_033_d2;
  assign _00070_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13505" *) _00641_ : vec_data_032_d2;
  assign _00068_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13495" *) _00640_ : vec_data_031_d2;
  assign _00066_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13485" *) _00639_ : vec_data_030_d2;
  assign _00064_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13475" *) _00638_ : vec_data_029_d2;
  assign _00062_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13465" *) _00637_ : vec_data_028_d2;
  assign _00060_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13455" *) _00636_ : vec_data_027_d2;
  assign _00058_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13445" *) _00635_ : vec_data_026_d2;
  assign _00056_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13435" *) _00634_ : vec_data_025_d2;
  assign _00054_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13425" *) _00633_ : vec_data_024_d2;
  assign _00052_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13415" *) _00632_ : vec_data_023_d2;
  assign _00050_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13405" *) _00631_ : vec_data_022_d2;
  assign _00048_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13395" *) _00630_ : vec_data_021_d2;
  assign _00046_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13385" *) _00629_ : vec_data_020_d2;
  assign _00044_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13375" *) _00628_ : vec_data_019_d2;
  assign _00042_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13365" *) _00627_ : vec_data_018_d2;
  assign _00040_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13355" *) _00626_ : vec_data_017_d2;
  assign _00038_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13345" *) _00625_ : vec_data_016_d2;
  assign _00036_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13335" *) _00624_ : vec_data_015_d2;
  assign _00034_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13325" *) _00623_ : vec_data_014_d2;
  assign _00032_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13315" *) _00622_ : vec_data_013_d2;
  assign _00030_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13305" *) _00621_ : vec_data_012_d2;
  assign _00028_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13295" *) _00620_ : vec_data_011_d2;
  assign _00026_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13285" *) _00619_ : vec_data_010_d2;
  assign _00024_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13275" *) _00618_ : vec_data_009_d2;
  assign _00022_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13265" *) _00617_ : vec_data_008_d2;
  assign _00020_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13255" *) _00616_ : vec_data_007_d2;
  assign _00018_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13245" *) _00615_ : vec_data_006_d2;
  assign _00016_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13235" *) _00614_ : vec_data_005_d2;
  assign _00014_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13225" *) _00613_ : vec_data_004_d2;
  assign _00012_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13215" *) _00612_ : vec_data_003_d2;
  assign _00010_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13205" *) _00611_ : vec_data_002_d2;
  assign _00008_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13195" *) _00610_ : vec_data_001_d2;
  assign _00006_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13185" *) _00609_ : vec_data_000_d2;
  assign _00004_ = valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13175" *) sel_d1 : sel_d2;
  function [7:0] _10136_;
    input [7:0] a;
    input [1023:0] b;
    input [127:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *)
    (* parallel_case *)
    casez (s)
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10136_ = b[7:0];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10136_ = b[15:8];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10136_ = b[23:16];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10136_ = b[31:24];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10136_ = b[39:32];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10136_ = b[47:40];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10136_ = b[55:48];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10136_ = b[63:56];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10136_ = b[71:64];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10136_ = b[79:72];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10136_ = b[87:80];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10136_ = b[95:88];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10136_ = b[103:96];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10136_ = b[111:104];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10136_ = b[119:112];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10136_ = b[127:120];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10136_ = b[135:128];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10136_ = b[143:136];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10136_ = b[151:144];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10136_ = b[159:152];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10136_ = b[167:160];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10136_ = b[175:168];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10136_ = b[183:176];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10136_ = b[191:184];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10136_ = b[199:192];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10136_ = b[207:200];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10136_ = b[215:208];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10136_ = b[223:216];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10136_ = b[231:224];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10136_ = b[239:232];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10136_ = b[247:240];
      128'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10136_ = b[255:248];
      128'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10136_ = b[263:256];
      128'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10136_ = b[271:264];
      128'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10136_ = b[279:272];
      128'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10136_ = b[287:280];
      128'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10136_ = b[295:288];
      128'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10136_ = b[303:296];
      128'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10136_ = b[311:304];
      128'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10136_ = b[319:312];
      128'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10136_ = b[327:320];
      128'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10136_ = b[335:328];
      128'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10136_ = b[343:336];
      128'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10136_ = b[351:344];
      128'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10136_ = b[359:352];
      128'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10136_ = b[367:360];
      128'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10136_ = b[375:368];
      128'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10136_ = b[383:376];
      128'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10136_ = b[391:384];
      128'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10136_ = b[399:392];
      128'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10136_ = b[407:400];
      128'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10136_ = b[415:408];
      128'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10136_ = b[423:416];
      128'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10136_ = b[431:424];
      128'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10136_ = b[439:432];
      128'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10136_ = b[447:440];
      128'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10136_ = b[455:448];
      128'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10136_ = b[463:456];
      128'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10136_ = b[471:464];
      128'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10136_ = b[479:472];
      128'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10136_ = b[487:480];
      128'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10136_ = b[495:488];
      128'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10136_ = b[503:496];
      128'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10136_ = b[511:504];
      128'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10136_ = b[519:512];
      128'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10136_ = b[527:520];
      128'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10136_ = b[535:528];
      128'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10136_ = b[543:536];
      128'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10136_ = b[551:544];
      128'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10136_ = b[559:552];
      128'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10136_ = b[567:560];
      128'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10136_ = b[575:568];
      128'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10136_ = b[583:576];
      128'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10136_ = b[591:584];
      128'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10136_ = b[599:592];
      128'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10136_ = b[607:600];
      128'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[615:608];
      128'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[623:616];
      128'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[631:624];
      128'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[639:632];
      128'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[647:640];
      128'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[655:648];
      128'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[663:656];
      128'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[671:664];
      128'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[679:672];
      128'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[687:680];
      128'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[695:688];
      128'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[703:696];
      128'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[711:704];
      128'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[719:712];
      128'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[727:720];
      128'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[735:728];
      128'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[743:736];
      128'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[751:744];
      128'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[759:752];
      128'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[767:760];
      128'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[775:768];
      128'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[783:776];
      128'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[791:784];
      128'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[799:792];
      128'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[807:800];
      128'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[815:808];
      128'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[823:816];
      128'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[831:824];
      128'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[839:832];
      128'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[847:840];
      128'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[855:848];
      128'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[863:856];
      128'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[871:864];
      128'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[879:872];
      128'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[887:880];
      128'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[895:888];
      128'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[903:896];
      128'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[911:904];
      128'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[919:912];
      128'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[927:920];
      128'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[935:928];
      128'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[943:936];
      128'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[951:944];
      128'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[959:952];
      128'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[967:960];
      128'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[975:968];
      128'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[983:976];
      128'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[991:984];
      128'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[999:992];
      128'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[1007:1000];
      128'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[1015:1008];
      128'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10136_ = b[1023:1016];
      default:
        _10136_ = a;
    endcase
  endfunction
  assign vec_data_127 = _10136_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976], data_d1[991:984], data_d1[999:992], data_d1[1007:1000], data_d1[1015:1008], data_d1[1023:1016] }, { _00873_, _00872_, _00871_, _00870_, _00869_, _00868_, _00867_, _00866_, _00865_, _00864_, _00863_, _00862_, _00861_, _00860_, _00859_, _00858_, _00857_, _00856_, _00855_, _00854_, _00853_, _00852_, _00851_, _00850_, _00849_, _00848_, _00847_, _00846_, _00845_, _00844_, _00843_, _00842_, _00841_, _00840_, _00839_, _00838_, _00837_, _00836_, _00835_, _00834_, _00833_, _00832_, _00831_, _00830_, _00829_, _00828_, _00827_, _00826_, _00825_, _00824_, _00823_, _00822_, _00821_, _00820_, _00819_, _00818_, _00817_, _00816_, _00815_, _00814_, _00813_, _00812_, _00811_, _00810_, _00809_, _00808_, _00807_, _00806_, _00805_, _00804_, _00803_, _00802_, _00801_, _00800_, _00799_, _00798_, _00797_, _00796_, _00795_, _00794_, _00793_, _00792_, _00791_, _00790_, _00789_, _00788_, _00787_, _00786_, _00785_, _00784_, _00783_, _00782_, _00781_, _00780_, _00779_, _00778_, _00777_, _00776_, _00775_, _00774_, _00773_, _00772_, _00771_, _00770_, _00769_, _00768_, _00767_, _00766_, _00765_, _00764_, _00763_, _00762_, _00761_, _00760_, _00759_, _00758_, _00757_, _00756_, _00755_, _00754_, _00753_, _00752_, _00751_, _00750_, _00749_, _00748_, _00747_, _00746_ });
  assign _00746_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 8'b10000000;
  assign _00747_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111111;
  assign _00748_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111110;
  assign _00749_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111101;
  assign _00750_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111100;
  assign _00751_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111011;
  assign _00752_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111010;
  assign _00753_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111001;
  assign _00754_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1111000;
  assign _00755_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110111;
  assign _00756_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110110;
  assign _00757_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110101;
  assign _00758_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110100;
  assign _00759_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110011;
  assign _00760_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110010;
  assign _00761_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110001;
  assign _00762_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1110000;
  assign _00763_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101111;
  assign _00764_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101110;
  assign _00765_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101101;
  assign _00766_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101100;
  assign _00767_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101011;
  assign _00768_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101010;
  assign _00769_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101001;
  assign _00770_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1101000;
  assign _00771_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100111;
  assign _00772_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100110;
  assign _00773_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100101;
  assign _00774_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100100;
  assign _00775_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100011;
  assign _00776_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100010;
  assign _00777_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100001;
  assign _00778_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1100000;
  assign _00779_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011111;
  assign _00780_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011110;
  assign _00781_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011101;
  assign _00782_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011100;
  assign _00783_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011011;
  assign _00784_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011010;
  assign _00785_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011001;
  assign _00786_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1011000;
  assign _00787_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010111;
  assign _00788_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010110;
  assign _00789_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010101;
  assign _00790_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010100;
  assign _00791_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010011;
  assign _00792_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010010;
  assign _00793_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010001;
  assign _00794_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1010000;
  assign _00795_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001111;
  assign _00796_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001110;
  assign _00797_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001101;
  assign _00798_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001100;
  assign _00799_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001011;
  assign _00800_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001010;
  assign _00801_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001001;
  assign _00802_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1001000;
  assign _00803_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000111;
  assign _00804_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000110;
  assign _00805_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000101;
  assign _00806_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000100;
  assign _00807_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000011;
  assign _00808_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000010;
  assign _00809_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000001;
  assign _00810_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 7'b1000000;
  assign _00811_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111111;
  assign _00812_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111110;
  assign _00813_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111101;
  assign _00814_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111100;
  assign _00815_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111011;
  assign _00816_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111010;
  assign _00817_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111001;
  assign _00818_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b111000;
  assign _00819_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110111;
  assign _00820_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110110;
  assign _00821_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110101;
  assign _00822_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110100;
  assign _00823_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110011;
  assign _00824_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110010;
  assign _00825_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110001;
  assign _00826_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b110000;
  assign _00827_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101111;
  assign _00828_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101110;
  assign _00829_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101101;
  assign _00830_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101100;
  assign _00831_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101011;
  assign _00832_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101010;
  assign _00833_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101001;
  assign _00834_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b101000;
  assign _00835_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100111;
  assign _00836_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100110;
  assign _00837_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100101;
  assign _00838_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100100;
  assign _00839_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100011;
  assign _00840_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100010;
  assign _00841_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100001;
  assign _00842_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 6'b100000;
  assign _00843_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11111;
  assign _00844_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11110;
  assign _00845_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11101;
  assign _00846_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11100;
  assign _00847_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11011;
  assign _00848_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11010;
  assign _00849_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11001;
  assign _00850_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b11000;
  assign _00851_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10111;
  assign _00852_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10110;
  assign _00853_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10101;
  assign _00854_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10100;
  assign _00855_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10011;
  assign _00856_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10010;
  assign _00857_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10001;
  assign _00858_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 5'b10000;
  assign _00859_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1111;
  assign _00860_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1110;
  assign _00861_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1101;
  assign _00862_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1100;
  assign _00863_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1011;
  assign _00864_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1010;
  assign _00865_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1001;
  assign _00866_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 4'b1000;
  assign _00867_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 3'b111;
  assign _00868_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 3'b110;
  assign _00869_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 3'b101;
  assign _00870_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 3'b100;
  assign _00871_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 2'b11;
  assign _00872_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 2'b10;
  assign _00873_ = { _00745_[7], vec_sum_127_d1 } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13035" *) 1'b1;
  function [7:0] _10265_;
    input [7:0] a;
    input [1015:0] b;
    input [126:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *)
    (* parallel_case *)
    casez (s)
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10265_ = b[7:0];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10265_ = b[15:8];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10265_ = b[23:16];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10265_ = b[31:24];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10265_ = b[39:32];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10265_ = b[47:40];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10265_ = b[55:48];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10265_ = b[63:56];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10265_ = b[71:64];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10265_ = b[79:72];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10265_ = b[87:80];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10265_ = b[95:88];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10265_ = b[103:96];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10265_ = b[111:104];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10265_ = b[119:112];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10265_ = b[127:120];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10265_ = b[135:128];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10265_ = b[143:136];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10265_ = b[151:144];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10265_ = b[159:152];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10265_ = b[167:160];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10265_ = b[175:168];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10265_ = b[183:176];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10265_ = b[191:184];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10265_ = b[199:192];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10265_ = b[207:200];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10265_ = b[215:208];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10265_ = b[223:216];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10265_ = b[231:224];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10265_ = b[239:232];
      127'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10265_ = b[247:240];
      127'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10265_ = b[255:248];
      127'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10265_ = b[263:256];
      127'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10265_ = b[271:264];
      127'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10265_ = b[279:272];
      127'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10265_ = b[287:280];
      127'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10265_ = b[295:288];
      127'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10265_ = b[303:296];
      127'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10265_ = b[311:304];
      127'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10265_ = b[319:312];
      127'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10265_ = b[327:320];
      127'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10265_ = b[335:328];
      127'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10265_ = b[343:336];
      127'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10265_ = b[351:344];
      127'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10265_ = b[359:352];
      127'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10265_ = b[367:360];
      127'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10265_ = b[375:368];
      127'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10265_ = b[383:376];
      127'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10265_ = b[391:384];
      127'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10265_ = b[399:392];
      127'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10265_ = b[407:400];
      127'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10265_ = b[415:408];
      127'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10265_ = b[423:416];
      127'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10265_ = b[431:424];
      127'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10265_ = b[439:432];
      127'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10265_ = b[447:440];
      127'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10265_ = b[455:448];
      127'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10265_ = b[463:456];
      127'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10265_ = b[471:464];
      127'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10265_ = b[479:472];
      127'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10265_ = b[487:480];
      127'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10265_ = b[495:488];
      127'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10265_ = b[503:496];
      127'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10265_ = b[511:504];
      127'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10265_ = b[519:512];
      127'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10265_ = b[527:520];
      127'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10265_ = b[535:528];
      127'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10265_ = b[543:536];
      127'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10265_ = b[551:544];
      127'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10265_ = b[559:552];
      127'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10265_ = b[567:560];
      127'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10265_ = b[575:568];
      127'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10265_ = b[583:576];
      127'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10265_ = b[591:584];
      127'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10265_ = b[599:592];
      127'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10265_ = b[607:600];
      127'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[615:608];
      127'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[623:616];
      127'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[631:624];
      127'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[639:632];
      127'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[647:640];
      127'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[655:648];
      127'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[663:656];
      127'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[671:664];
      127'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[679:672];
      127'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[687:680];
      127'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[695:688];
      127'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[703:696];
      127'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[711:704];
      127'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[719:712];
      127'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[727:720];
      127'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[735:728];
      127'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[743:736];
      127'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[751:744];
      127'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[759:752];
      127'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[767:760];
      127'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[775:768];
      127'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[783:776];
      127'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[791:784];
      127'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[799:792];
      127'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[807:800];
      127'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[815:808];
      127'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[823:816];
      127'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[831:824];
      127'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[839:832];
      127'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[847:840];
      127'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[855:848];
      127'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[863:856];
      127'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[871:864];
      127'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[879:872];
      127'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[887:880];
      127'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[895:888];
      127'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[903:896];
      127'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[911:904];
      127'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[919:912];
      127'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[927:920];
      127'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[935:928];
      127'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[943:936];
      127'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[951:944];
      127'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[959:952];
      127'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[967:960];
      127'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[975:968];
      127'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[983:976];
      127'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[991:984];
      127'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[999:992];
      127'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[1007:1000];
      127'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10265_ = b[1015:1008];
      default:
        _10265_ = a;
    endcase
  endfunction
  assign vec_data_126 = _10265_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976], data_d1[991:984], data_d1[999:992], data_d1[1007:1000], data_d1[1015:1008] }, { _01000_, _00999_, _00998_, _00997_, _00996_, _00995_, _00994_, _00993_, _00992_, _00991_, _00990_, _00989_, _00988_, _00987_, _00986_, _00985_, _00984_, _00983_, _00982_, _00981_, _00980_, _00979_, _00978_, _00977_, _00976_, _00975_, _00974_, _00973_, _00972_, _00971_, _00970_, _00969_, _00968_, _00967_, _00966_, _00965_, _00964_, _00963_, _00962_, _00961_, _00960_, _00959_, _00958_, _00957_, _00956_, _00955_, _00954_, _00953_, _00952_, _00951_, _00950_, _00949_, _00948_, _00947_, _00946_, _00945_, _00944_, _00943_, _00942_, _00941_, _00940_, _00939_, _00938_, _00937_, _00936_, _00935_, _00934_, _00933_, _00932_, _00931_, _00930_, _00929_, _00928_, _00927_, _00926_, _00925_, _00924_, _00923_, _00922_, _00921_, _00920_, _00919_, _00918_, _00917_, _00916_, _00915_, _00914_, _00913_, _00912_, _00911_, _00910_, _00909_, _00908_, _00907_, _00906_, _00905_, _00904_, _00903_, _00902_, _00901_, _00900_, _00899_, _00898_, _00897_, _00896_, _00895_, _00894_, _00893_, _00892_, _00891_, _00890_, _00889_, _00888_, _00887_, _00886_, _00885_, _00884_, _00883_, _00882_, _00881_, _00880_, _00879_, _00878_, _00877_, _00876_, _00875_, _00874_ });
  assign _00874_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111111;
  assign _00875_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111110;
  assign _00876_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111101;
  assign _00877_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111100;
  assign _00878_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111011;
  assign _00879_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111010;
  assign _00880_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111001;
  assign _00881_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1111000;
  assign _00882_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110111;
  assign _00883_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110110;
  assign _00884_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110101;
  assign _00885_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110100;
  assign _00886_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110011;
  assign _00887_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110010;
  assign _00888_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110001;
  assign _00889_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1110000;
  assign _00890_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101111;
  assign _00891_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101110;
  assign _00892_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101101;
  assign _00893_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101100;
  assign _00894_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101011;
  assign _00895_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101010;
  assign _00896_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101001;
  assign _00897_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1101000;
  assign _00898_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100111;
  assign _00899_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100110;
  assign _00900_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100101;
  assign _00901_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:13000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100100;
  assign _00902_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100011;
  assign _00903_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100010;
  assign _00904_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100001;
  assign _00905_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1100000;
  assign _00906_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011111;
  assign _00907_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011110;
  assign _00908_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011101;
  assign _00909_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011100;
  assign _00910_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011011;
  assign _00911_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011010;
  assign _00912_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011001;
  assign _00913_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1011000;
  assign _00914_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010111;
  assign _00915_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010110;
  assign _00916_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010101;
  assign _00917_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010100;
  assign _00918_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010011;
  assign _00919_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010010;
  assign _00920_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010001;
  assign _00921_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1010000;
  assign _00922_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001111;
  assign _00923_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001110;
  assign _00924_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001101;
  assign _00925_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001100;
  assign _00926_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001011;
  assign _00927_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001010;
  assign _00928_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001001;
  assign _00929_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1001000;
  assign _00930_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000111;
  assign _00931_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000110;
  assign _00932_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000101;
  assign _00933_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000100;
  assign _00934_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000011;
  assign _00935_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000010;
  assign _00936_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000001;
  assign _00937_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 7'b1000000;
  assign _00938_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111111;
  assign _00939_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111110;
  assign _00940_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111101;
  assign _00941_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111100;
  assign _00942_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111011;
  assign _00943_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111010;
  assign _00944_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111001;
  assign _00945_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b111000;
  assign _00946_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110111;
  assign _00947_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110110;
  assign _00948_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110101;
  assign _00949_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110100;
  assign _00950_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110011;
  assign _00951_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110010;
  assign _00952_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110001;
  assign _00953_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b110000;
  assign _00954_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101111;
  assign _00955_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101110;
  assign _00956_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101101;
  assign _00957_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101100;
  assign _00958_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101011;
  assign _00959_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101010;
  assign _00960_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101001;
  assign _00961_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b101000;
  assign _00962_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100111;
  assign _00963_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100110;
  assign _00964_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100101;
  assign _00965_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100100;
  assign _00966_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100011;
  assign _00967_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100010;
  assign _00968_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100001;
  assign _00969_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 6'b100000;
  assign _00970_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11111;
  assign _00971_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11110;
  assign _00972_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11101;
  assign _00973_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11100;
  assign _00974_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11011;
  assign _00975_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11010;
  assign _00976_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11001;
  assign _00977_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b11000;
  assign _00978_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10111;
  assign _00979_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10110;
  assign _00980_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10101;
  assign _00981_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10100;
  assign _00982_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10011;
  assign _00983_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10010;
  assign _00984_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10001;
  assign _00985_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 5'b10000;
  assign _00986_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1111;
  assign _00987_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1110;
  assign _00988_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1101;
  assign _00989_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1100;
  assign _00990_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1011;
  assign _00991_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1010;
  assign _00992_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1001;
  assign _00993_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 4'b1000;
  assign _00994_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 3'b111;
  assign _00995_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 3'b110;
  assign _00996_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 3'b101;
  assign _00997_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 3'b100;
  assign _00998_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 2'b11;
  assign _00999_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 2'b10;
  assign _01000_ = vec_sum_126_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12900" *) 1'b1;
  function [7:0] _10393_;
    input [7:0] a;
    input [1007:0] b;
    input [125:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *)
    (* parallel_case *)
    casez (s)
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10393_ = b[7:0];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10393_ = b[15:8];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10393_ = b[23:16];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10393_ = b[31:24];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10393_ = b[39:32];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10393_ = b[47:40];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10393_ = b[55:48];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10393_ = b[63:56];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10393_ = b[71:64];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10393_ = b[79:72];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10393_ = b[87:80];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10393_ = b[95:88];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10393_ = b[103:96];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10393_ = b[111:104];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10393_ = b[119:112];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10393_ = b[127:120];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10393_ = b[135:128];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10393_ = b[143:136];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10393_ = b[151:144];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10393_ = b[159:152];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10393_ = b[167:160];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10393_ = b[175:168];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10393_ = b[183:176];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10393_ = b[191:184];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10393_ = b[199:192];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10393_ = b[207:200];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10393_ = b[215:208];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10393_ = b[223:216];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10393_ = b[231:224];
      126'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10393_ = b[239:232];
      126'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10393_ = b[247:240];
      126'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10393_ = b[255:248];
      126'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10393_ = b[263:256];
      126'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10393_ = b[271:264];
      126'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10393_ = b[279:272];
      126'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10393_ = b[287:280];
      126'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10393_ = b[295:288];
      126'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10393_ = b[303:296];
      126'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10393_ = b[311:304];
      126'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10393_ = b[319:312];
      126'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10393_ = b[327:320];
      126'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10393_ = b[335:328];
      126'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10393_ = b[343:336];
      126'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10393_ = b[351:344];
      126'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10393_ = b[359:352];
      126'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10393_ = b[367:360];
      126'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10393_ = b[375:368];
      126'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10393_ = b[383:376];
      126'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10393_ = b[391:384];
      126'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10393_ = b[399:392];
      126'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10393_ = b[407:400];
      126'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10393_ = b[415:408];
      126'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10393_ = b[423:416];
      126'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10393_ = b[431:424];
      126'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10393_ = b[439:432];
      126'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10393_ = b[447:440];
      126'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10393_ = b[455:448];
      126'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10393_ = b[463:456];
      126'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10393_ = b[471:464];
      126'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10393_ = b[479:472];
      126'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10393_ = b[487:480];
      126'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10393_ = b[495:488];
      126'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10393_ = b[503:496];
      126'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10393_ = b[511:504];
      126'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10393_ = b[519:512];
      126'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10393_ = b[527:520];
      126'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10393_ = b[535:528];
      126'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10393_ = b[543:536];
      126'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10393_ = b[551:544];
      126'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10393_ = b[559:552];
      126'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10393_ = b[567:560];
      126'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10393_ = b[575:568];
      126'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10393_ = b[583:576];
      126'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10393_ = b[591:584];
      126'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10393_ = b[599:592];
      126'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10393_ = b[607:600];
      126'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[615:608];
      126'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[623:616];
      126'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[631:624];
      126'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[639:632];
      126'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[647:640];
      126'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[655:648];
      126'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[663:656];
      126'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[671:664];
      126'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[679:672];
      126'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[687:680];
      126'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[695:688];
      126'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[703:696];
      126'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[711:704];
      126'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[719:712];
      126'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[727:720];
      126'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[735:728];
      126'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[743:736];
      126'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[751:744];
      126'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[759:752];
      126'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[767:760];
      126'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[775:768];
      126'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[783:776];
      126'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[791:784];
      126'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[799:792];
      126'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[807:800];
      126'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[815:808];
      126'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[823:816];
      126'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[831:824];
      126'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[839:832];
      126'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[847:840];
      126'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[855:848];
      126'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[863:856];
      126'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[871:864];
      126'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[879:872];
      126'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[887:880];
      126'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[895:888];
      126'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[903:896];
      126'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[911:904];
      126'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[919:912];
      126'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[927:920];
      126'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[935:928];
      126'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[943:936];
      126'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[951:944];
      126'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[959:952];
      126'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[967:960];
      126'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[975:968];
      126'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[983:976];
      126'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[991:984];
      126'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[999:992];
      126'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10393_ = b[1007:1000];
      default:
        _10393_ = a;
    endcase
  endfunction
  assign vec_data_125 = _10393_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976], data_d1[991:984], data_d1[999:992], data_d1[1007:1000] }, { _01126_, _01125_, _01124_, _01123_, _01122_, _01121_, _01120_, _01119_, _01118_, _01117_, _01116_, _01115_, _01114_, _01113_, _01112_, _01111_, _01110_, _01109_, _01108_, _01107_, _01106_, _01105_, _01104_, _01103_, _01102_, _01101_, _01100_, _01099_, _01098_, _01097_, _01096_, _01095_, _01094_, _01093_, _01092_, _01091_, _01090_, _01089_, _01088_, _01087_, _01086_, _01085_, _01084_, _01083_, _01082_, _01081_, _01080_, _01079_, _01078_, _01077_, _01076_, _01075_, _01074_, _01073_, _01072_, _01071_, _01070_, _01069_, _01068_, _01067_, _01066_, _01065_, _01064_, _01063_, _01062_, _01061_, _01060_, _01059_, _01058_, _01057_, _01056_, _01055_, _01054_, _01053_, _01052_, _01051_, _01050_, _01049_, _01048_, _01047_, _01046_, _01045_, _01044_, _01043_, _01042_, _01041_, _01040_, _01039_, _01038_, _01037_, _01036_, _01035_, _01034_, _01033_, _01032_, _01031_, _01030_, _01029_, _01028_, _01027_, _01026_, _01025_, _01024_, _01023_, _01022_, _01021_, _01020_, _01019_, _01018_, _01017_, _01016_, _01015_, _01014_, _01013_, _01012_, _01011_, _01010_, _01009_, _01008_, _01007_, _01006_, _01005_, _01004_, _01003_, _01002_, _01001_ });
  assign _01001_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111110;
  assign _01002_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111101;
  assign _01003_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111100;
  assign _01004_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111011;
  assign _01005_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111010;
  assign _01006_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111001;
  assign _01007_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1111000;
  assign _01008_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110111;
  assign _01009_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110110;
  assign _01010_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110101;
  assign _01011_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110100;
  assign _01012_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110011;
  assign _01013_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110010;
  assign _01014_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110001;
  assign _01015_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1110000;
  assign _01016_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101111;
  assign _01017_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101110;
  assign _01018_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101101;
  assign _01019_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101100;
  assign _01020_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101011;
  assign _01021_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101010;
  assign _01022_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101001;
  assign _01023_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1101000;
  assign _01024_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100111;
  assign _01025_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100110;
  assign _01026_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100101;
  assign _01027_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100100;
  assign _01028_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100011;
  assign _01029_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100010;
  assign _01030_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100001;
  assign _01031_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1100000;
  assign _01032_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011111;
  assign _01033_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011110;
  assign _01034_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011101;
  assign _01035_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011100;
  assign _01036_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011011;
  assign _01037_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011010;
  assign _01038_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011001;
  assign _01039_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1011000;
  assign _01040_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010111;
  assign _01041_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010110;
  assign _01042_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010101;
  assign _01043_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010100;
  assign _01044_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010011;
  assign _01045_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010010;
  assign _01046_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010001;
  assign _01047_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1010000;
  assign _01048_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001111;
  assign _01049_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001110;
  assign _01050_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001101;
  assign _01051_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001100;
  assign _01052_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001011;
  assign _01053_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001010;
  assign _01054_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001001;
  assign _01055_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1001000;
  assign _01056_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000111;
  assign _01057_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000110;
  assign _01058_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000101;
  assign _01059_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000100;
  assign _01060_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000011;
  assign _01061_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000010;
  assign _01062_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000001;
  assign _01063_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 7'b1000000;
  assign _01064_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111111;
  assign _01065_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111110;
  assign _01066_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111101;
  assign _01067_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111100;
  assign _01068_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111011;
  assign _01069_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111010;
  assign _01070_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111001;
  assign _01071_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b111000;
  assign _01072_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110111;
  assign _01073_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110110;
  assign _01074_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110101;
  assign _01075_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110100;
  assign _01076_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110011;
  assign _01077_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110010;
  assign _01078_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110001;
  assign _01079_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b110000;
  assign _01080_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101111;
  assign _01081_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101110;
  assign _01082_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101101;
  assign _01083_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101100;
  assign _01084_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101011;
  assign _01085_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101010;
  assign _01086_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101001;
  assign _01087_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b101000;
  assign _01088_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100111;
  assign _01089_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100110;
  assign _01090_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100101;
  assign _01091_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100100;
  assign _01092_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100011;
  assign _01093_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100010;
  assign _01094_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100001;
  assign _01095_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 6'b100000;
  assign _01096_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11111;
  assign _01097_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11110;
  assign _01098_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11101;
  assign _01099_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11100;
  assign _01100_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11011;
  assign _01101_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11010;
  assign _01102_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11001;
  assign _01103_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b11000;
  assign _01104_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10111;
  assign _01105_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10110;
  assign _01106_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10101;
  assign _01107_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10100;
  assign _01108_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10011;
  assign _01109_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10010;
  assign _01110_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10001;
  assign _01111_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 5'b10000;
  assign _01112_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1111;
  assign _01113_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1110;
  assign _01114_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1101;
  assign _01115_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1100;
  assign _01116_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1011;
  assign _01117_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1010;
  assign _01118_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1001;
  assign _01119_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 4'b1000;
  assign _01120_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 3'b111;
  assign _01121_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 3'b110;
  assign _01122_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 3'b101;
  assign _01123_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 3'b100;
  assign _01124_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 2'b11;
  assign _01125_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 2'b10;
  assign _01126_ = vec_sum_125_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12766" *) 1'b1;
  function [7:0] _10520_;
    input [7:0] a;
    input [999:0] b;
    input [124:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *)
    (* parallel_case *)
    casez (s)
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10520_ = b[7:0];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10520_ = b[15:8];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10520_ = b[23:16];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10520_ = b[31:24];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10520_ = b[39:32];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10520_ = b[47:40];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10520_ = b[55:48];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10520_ = b[63:56];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10520_ = b[71:64];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10520_ = b[79:72];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10520_ = b[87:80];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10520_ = b[95:88];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10520_ = b[103:96];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10520_ = b[111:104];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10520_ = b[119:112];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10520_ = b[127:120];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10520_ = b[135:128];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10520_ = b[143:136];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10520_ = b[151:144];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10520_ = b[159:152];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10520_ = b[167:160];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10520_ = b[175:168];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10520_ = b[183:176];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10520_ = b[191:184];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10520_ = b[199:192];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10520_ = b[207:200];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10520_ = b[215:208];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10520_ = b[223:216];
      125'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10520_ = b[231:224];
      125'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10520_ = b[239:232];
      125'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10520_ = b[247:240];
      125'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10520_ = b[255:248];
      125'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10520_ = b[263:256];
      125'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10520_ = b[271:264];
      125'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10520_ = b[279:272];
      125'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10520_ = b[287:280];
      125'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10520_ = b[295:288];
      125'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10520_ = b[303:296];
      125'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10520_ = b[311:304];
      125'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10520_ = b[319:312];
      125'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10520_ = b[327:320];
      125'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10520_ = b[335:328];
      125'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10520_ = b[343:336];
      125'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10520_ = b[351:344];
      125'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10520_ = b[359:352];
      125'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10520_ = b[367:360];
      125'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10520_ = b[375:368];
      125'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10520_ = b[383:376];
      125'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10520_ = b[391:384];
      125'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10520_ = b[399:392];
      125'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10520_ = b[407:400];
      125'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10520_ = b[415:408];
      125'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10520_ = b[423:416];
      125'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10520_ = b[431:424];
      125'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10520_ = b[439:432];
      125'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10520_ = b[447:440];
      125'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10520_ = b[455:448];
      125'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10520_ = b[463:456];
      125'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10520_ = b[471:464];
      125'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10520_ = b[479:472];
      125'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10520_ = b[487:480];
      125'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10520_ = b[495:488];
      125'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10520_ = b[503:496];
      125'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10520_ = b[511:504];
      125'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10520_ = b[519:512];
      125'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10520_ = b[527:520];
      125'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10520_ = b[535:528];
      125'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10520_ = b[543:536];
      125'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10520_ = b[551:544];
      125'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10520_ = b[559:552];
      125'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10520_ = b[567:560];
      125'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10520_ = b[575:568];
      125'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10520_ = b[583:576];
      125'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10520_ = b[591:584];
      125'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10520_ = b[599:592];
      125'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10520_ = b[607:600];
      125'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[615:608];
      125'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[623:616];
      125'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[631:624];
      125'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[639:632];
      125'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[647:640];
      125'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[655:648];
      125'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[663:656];
      125'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[671:664];
      125'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[679:672];
      125'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[687:680];
      125'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[695:688];
      125'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[703:696];
      125'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[711:704];
      125'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[719:712];
      125'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[727:720];
      125'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[735:728];
      125'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[743:736];
      125'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[751:744];
      125'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[759:752];
      125'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[767:760];
      125'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[775:768];
      125'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[783:776];
      125'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[791:784];
      125'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[799:792];
      125'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[807:800];
      125'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[815:808];
      125'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[823:816];
      125'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[831:824];
      125'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[839:832];
      125'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[847:840];
      125'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[855:848];
      125'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[863:856];
      125'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[871:864];
      125'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[879:872];
      125'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[887:880];
      125'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[895:888];
      125'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[903:896];
      125'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[911:904];
      125'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[919:912];
      125'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[927:920];
      125'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[935:928];
      125'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[943:936];
      125'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[951:944];
      125'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[959:952];
      125'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[967:960];
      125'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[975:968];
      125'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[983:976];
      125'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[991:984];
      125'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10520_ = b[999:992];
      default:
        _10520_ = a;
    endcase
  endfunction
  assign vec_data_124 = _10520_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976], data_d1[991:984], data_d1[999:992] }, { _01251_, _01250_, _01249_, _01248_, _01247_, _01246_, _01245_, _01244_, _01243_, _01242_, _01241_, _01240_, _01239_, _01238_, _01237_, _01236_, _01235_, _01234_, _01233_, _01232_, _01231_, _01230_, _01229_, _01228_, _01227_, _01226_, _01225_, _01224_, _01223_, _01222_, _01221_, _01220_, _01219_, _01218_, _01217_, _01216_, _01215_, _01214_, _01213_, _01212_, _01211_, _01210_, _01209_, _01208_, _01207_, _01206_, _01205_, _01204_, _01203_, _01202_, _01201_, _01200_, _01199_, _01198_, _01197_, _01196_, _01195_, _01194_, _01193_, _01192_, _01191_, _01190_, _01189_, _01188_, _01187_, _01186_, _01185_, _01184_, _01183_, _01182_, _01181_, _01180_, _01179_, _01178_, _01177_, _01176_, _01175_, _01174_, _01173_, _01172_, _01171_, _01170_, _01169_, _01168_, _01167_, _01166_, _01165_, _01164_, _01163_, _01162_, _01161_, _01160_, _01159_, _01158_, _01157_, _01156_, _01155_, _01154_, _01153_, _01152_, _01151_, _01150_, _01149_, _01148_, _01147_, _01146_, _01145_, _01144_, _01143_, _01142_, _01141_, _01140_, _01139_, _01138_, _01137_, _01136_, _01135_, _01134_, _01133_, _01132_, _01131_, _01130_, _01129_, _01128_, _01127_ });
  assign _01127_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111101;
  assign _01128_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111100;
  assign _01129_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111011;
  assign _01130_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111010;
  assign _01131_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111001;
  assign _01132_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1111000;
  assign _01133_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110111;
  assign _01134_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110110;
  assign _01135_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110101;
  assign _01136_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110100;
  assign _01137_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110011;
  assign _01138_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110010;
  assign _01139_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110001;
  assign _01140_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1110000;
  assign _01141_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101111;
  assign _01142_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101110;
  assign _01143_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101101;
  assign _01144_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101100;
  assign _01145_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101011;
  assign _01146_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101010;
  assign _01147_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101001;
  assign _01148_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1101000;
  assign _01149_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100111;
  assign _01150_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100110;
  assign _01151_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100101;
  assign _01152_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100100;
  assign _01153_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100011;
  assign _01154_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100010;
  assign _01155_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100001;
  assign _01156_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1100000;
  assign _01157_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011111;
  assign _01158_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011110;
  assign _01159_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011101;
  assign _01160_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011100;
  assign _01161_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011011;
  assign _01162_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011010;
  assign _01163_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011001;
  assign _01164_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1011000;
  assign _01165_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010111;
  assign _01166_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010110;
  assign _01167_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010101;
  assign _01168_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010100;
  assign _01169_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010011;
  assign _01170_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010010;
  assign _01171_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010001;
  assign _01172_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1010000;
  assign _01173_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001111;
  assign _01174_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001110;
  assign _01175_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001101;
  assign _01176_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001100;
  assign _01177_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001011;
  assign _01178_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001010;
  assign _01179_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001001;
  assign _01180_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1001000;
  assign _01181_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000111;
  assign _01182_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000110;
  assign _01183_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000101;
  assign _01184_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000100;
  assign _01185_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000011;
  assign _01186_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000010;
  assign _01187_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000001;
  assign _01188_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 7'b1000000;
  assign _01189_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111111;
  assign _01190_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111110;
  assign _01191_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111101;
  assign _01192_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111100;
  assign _01193_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111011;
  assign _01194_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111010;
  assign _01195_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111001;
  assign _01196_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b111000;
  assign _01197_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110111;
  assign _01198_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110110;
  assign _01199_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110101;
  assign _01200_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110100;
  assign _01201_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110011;
  assign _01202_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110010;
  assign _01203_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110001;
  assign _01204_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b110000;
  assign _01205_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101111;
  assign _01206_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101110;
  assign _01207_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101101;
  assign _01208_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101100;
  assign _01209_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101011;
  assign _01210_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101010;
  assign _01211_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101001;
  assign _01212_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b101000;
  assign _01213_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100111;
  assign _01214_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100110;
  assign _01215_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100101;
  assign _01216_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100100;
  assign _01217_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100011;
  assign _01218_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100010;
  assign _01219_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100001;
  assign _01220_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 6'b100000;
  assign _01221_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11111;
  assign _01222_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11110;
  assign _01223_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11101;
  assign _01224_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11100;
  assign _01225_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11011;
  assign _01226_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11010;
  assign _01227_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11001;
  assign _01228_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b11000;
  assign _01229_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10111;
  assign _01230_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10110;
  assign _01231_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10101;
  assign _01232_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10100;
  assign _01233_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10011;
  assign _01234_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10010;
  assign _01235_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10001;
  assign _01236_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 5'b10000;
  assign _01237_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1111;
  assign _01238_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1110;
  assign _01239_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1101;
  assign _01240_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1100;
  assign _01241_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1011;
  assign _01242_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1010;
  assign _01243_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1001;
  assign _01244_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 4'b1000;
  assign _01245_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 3'b111;
  assign _01246_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 3'b110;
  assign _01247_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 3'b101;
  assign _01248_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 3'b100;
  assign _01249_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 2'b11;
  assign _01250_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 2'b10;
  assign _01251_ = vec_sum_124_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12633" *) 1'b1;
  function [7:0] _10646_;
    input [7:0] a;
    input [991:0] b;
    input [123:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *)
    (* parallel_case *)
    casez (s)
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10646_ = b[7:0];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10646_ = b[15:8];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10646_ = b[23:16];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10646_ = b[31:24];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10646_ = b[39:32];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10646_ = b[47:40];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10646_ = b[55:48];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10646_ = b[63:56];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10646_ = b[71:64];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10646_ = b[79:72];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10646_ = b[87:80];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10646_ = b[95:88];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10646_ = b[103:96];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10646_ = b[111:104];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10646_ = b[119:112];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10646_ = b[127:120];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10646_ = b[135:128];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10646_ = b[143:136];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10646_ = b[151:144];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10646_ = b[159:152];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10646_ = b[167:160];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10646_ = b[175:168];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10646_ = b[183:176];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10646_ = b[191:184];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10646_ = b[199:192];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10646_ = b[207:200];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10646_ = b[215:208];
      124'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10646_ = b[223:216];
      124'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10646_ = b[231:224];
      124'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10646_ = b[239:232];
      124'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10646_ = b[247:240];
      124'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10646_ = b[255:248];
      124'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10646_ = b[263:256];
      124'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10646_ = b[271:264];
      124'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10646_ = b[279:272];
      124'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10646_ = b[287:280];
      124'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10646_ = b[295:288];
      124'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10646_ = b[303:296];
      124'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10646_ = b[311:304];
      124'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10646_ = b[319:312];
      124'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10646_ = b[327:320];
      124'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10646_ = b[335:328];
      124'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10646_ = b[343:336];
      124'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10646_ = b[351:344];
      124'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10646_ = b[359:352];
      124'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10646_ = b[367:360];
      124'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10646_ = b[375:368];
      124'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10646_ = b[383:376];
      124'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10646_ = b[391:384];
      124'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10646_ = b[399:392];
      124'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10646_ = b[407:400];
      124'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10646_ = b[415:408];
      124'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10646_ = b[423:416];
      124'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10646_ = b[431:424];
      124'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10646_ = b[439:432];
      124'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10646_ = b[447:440];
      124'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10646_ = b[455:448];
      124'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10646_ = b[463:456];
      124'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10646_ = b[471:464];
      124'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10646_ = b[479:472];
      124'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10646_ = b[487:480];
      124'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10646_ = b[495:488];
      124'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10646_ = b[503:496];
      124'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10646_ = b[511:504];
      124'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10646_ = b[519:512];
      124'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10646_ = b[527:520];
      124'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10646_ = b[535:528];
      124'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10646_ = b[543:536];
      124'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10646_ = b[551:544];
      124'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10646_ = b[559:552];
      124'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10646_ = b[567:560];
      124'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10646_ = b[575:568];
      124'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10646_ = b[583:576];
      124'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10646_ = b[591:584];
      124'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10646_ = b[599:592];
      124'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10646_ = b[607:600];
      124'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[615:608];
      124'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[623:616];
      124'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[631:624];
      124'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[639:632];
      124'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[647:640];
      124'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[655:648];
      124'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[663:656];
      124'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[671:664];
      124'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[679:672];
      124'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[687:680];
      124'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[695:688];
      124'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[703:696];
      124'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[711:704];
      124'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[719:712];
      124'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[727:720];
      124'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[735:728];
      124'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[743:736];
      124'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[751:744];
      124'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[759:752];
      124'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[767:760];
      124'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[775:768];
      124'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[783:776];
      124'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[791:784];
      124'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[799:792];
      124'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[807:800];
      124'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[815:808];
      124'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[823:816];
      124'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[831:824];
      124'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[839:832];
      124'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[847:840];
      124'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[855:848];
      124'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[863:856];
      124'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[871:864];
      124'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[879:872];
      124'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[887:880];
      124'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[895:888];
      124'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[903:896];
      124'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[911:904];
      124'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[919:912];
      124'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[927:920];
      124'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[935:928];
      124'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[943:936];
      124'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[951:944];
      124'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[959:952];
      124'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[967:960];
      124'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[975:968];
      124'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[983:976];
      124'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10646_ = b[991:984];
      default:
        _10646_ = a;
    endcase
  endfunction
  assign vec_data_123 = _10646_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976], data_d1[991:984] }, { _01375_, _01374_, _01373_, _01372_, _01371_, _01370_, _01369_, _01368_, _01367_, _01366_, _01365_, _01364_, _01363_, _01362_, _01361_, _01360_, _01359_, _01358_, _01357_, _01356_, _01355_, _01354_, _01353_, _01352_, _01351_, _01350_, _01349_, _01348_, _01347_, _01346_, _01345_, _01344_, _01343_, _01342_, _01341_, _01340_, _01339_, _01338_, _01337_, _01336_, _01335_, _01334_, _01333_, _01332_, _01331_, _01330_, _01329_, _01328_, _01327_, _01326_, _01325_, _01324_, _01323_, _01322_, _01321_, _01320_, _01319_, _01318_, _01317_, _01316_, _01315_, _01314_, _01313_, _01312_, _01311_, _01310_, _01309_, _01308_, _01307_, _01306_, _01305_, _01304_, _01303_, _01302_, _01301_, _01300_, _01299_, _01298_, _01297_, _01296_, _01295_, _01294_, _01293_, _01292_, _01291_, _01290_, _01289_, _01288_, _01287_, _01286_, _01285_, _01284_, _01283_, _01282_, _01281_, _01280_, _01279_, _01278_, _01277_, _01276_, _01275_, _01274_, _01273_, _01272_, _01271_, _01270_, _01269_, _01268_, _01267_, _01266_, _01265_, _01264_, _01263_, _01262_, _01261_, _01260_, _01259_, _01258_, _01257_, _01256_, _01255_, _01254_, _01253_, _01252_ });
  assign _01252_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1111100;
  assign _01253_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1111011;
  assign _01254_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1111010;
  assign _01255_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1111001;
  assign _01256_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1111000;
  assign _01257_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110111;
  assign _01258_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110110;
  assign _01259_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110101;
  assign _01260_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110100;
  assign _01261_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110011;
  assign _01262_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110010;
  assign _01263_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110001;
  assign _01264_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1110000;
  assign _01265_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101111;
  assign _01266_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101110;
  assign _01267_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101101;
  assign _01268_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101100;
  assign _01269_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101011;
  assign _01270_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101010;
  assign _01271_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101001;
  assign _01272_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1101000;
  assign _01273_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100111;
  assign _01274_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100110;
  assign _01275_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100101;
  assign _01276_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100100;
  assign _01277_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100011;
  assign _01278_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100010;
  assign _01279_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100001;
  assign _01280_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1100000;
  assign _01281_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011111;
  assign _01282_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011110;
  assign _01283_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011101;
  assign _01284_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011100;
  assign _01285_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011011;
  assign _01286_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011010;
  assign _01287_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011001;
  assign _01288_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1011000;
  assign _01289_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010111;
  assign _01290_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010110;
  assign _01291_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010101;
  assign _01292_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010100;
  assign _01293_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010011;
  assign _01294_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010010;
  assign _01295_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010001;
  assign _01296_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1010000;
  assign _01297_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001111;
  assign _01298_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001110;
  assign _01299_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001101;
  assign _01300_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001100;
  assign _01301_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001011;
  assign _01302_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001010;
  assign _01303_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001001;
  assign _01304_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1001000;
  assign _01305_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000111;
  assign _01306_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000110;
  assign _01307_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000101;
  assign _01308_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000100;
  assign _01309_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000011;
  assign _01310_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000010;
  assign _01311_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000001;
  assign _01312_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 7'b1000000;
  assign _01313_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111111;
  assign _01314_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111110;
  assign _01315_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111101;
  assign _01316_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111100;
  assign _01317_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111011;
  assign _01318_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111010;
  assign _01319_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111001;
  assign _01320_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b111000;
  assign _01321_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110111;
  assign _01322_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110110;
  assign _01323_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110101;
  assign _01324_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110100;
  assign _01325_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110011;
  assign _01326_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110010;
  assign _01327_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110001;
  assign _01328_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b110000;
  assign _01329_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101111;
  assign _01330_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101110;
  assign _01331_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101101;
  assign _01332_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101100;
  assign _01333_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101011;
  assign _01334_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101010;
  assign _01335_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101001;
  assign _01336_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b101000;
  assign _01337_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100111;
  assign _01338_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100110;
  assign _01339_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100101;
  assign _01340_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100100;
  assign _01341_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100011;
  assign _01342_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100010;
  assign _01343_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100001;
  assign _01344_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 6'b100000;
  assign _01345_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11111;
  assign _01346_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11110;
  assign _01347_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11101;
  assign _01348_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11100;
  assign _01349_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11011;
  assign _01350_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11010;
  assign _01351_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11001;
  assign _01352_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b11000;
  assign _01353_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10111;
  assign _01354_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10110;
  assign _01355_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10101;
  assign _01356_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10100;
  assign _01357_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10011;
  assign _01358_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10010;
  assign _01359_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10001;
  assign _01360_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 5'b10000;
  assign _01361_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1111;
  assign _01362_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1110;
  assign _01363_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1101;
  assign _01364_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1100;
  assign _01365_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1011;
  assign _01366_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1010;
  assign _01367_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1001;
  assign _01368_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 4'b1000;
  assign _01369_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 3'b111;
  assign _01370_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 3'b110;
  assign _01371_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 3'b101;
  assign _01372_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 3'b100;
  assign _01373_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 2'b11;
  assign _01374_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 2'b10;
  assign _01375_ = vec_sum_123_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12501" *) 1'b1;
  function [7:0] _10771_;
    input [7:0] a;
    input [983:0] b;
    input [122:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *)
    (* parallel_case *)
    casez (s)
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10771_ = b[7:0];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10771_ = b[15:8];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10771_ = b[23:16];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10771_ = b[31:24];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10771_ = b[39:32];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10771_ = b[47:40];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10771_ = b[55:48];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10771_ = b[63:56];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10771_ = b[71:64];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10771_ = b[79:72];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10771_ = b[87:80];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10771_ = b[95:88];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10771_ = b[103:96];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10771_ = b[111:104];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10771_ = b[119:112];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10771_ = b[127:120];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10771_ = b[135:128];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10771_ = b[143:136];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10771_ = b[151:144];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10771_ = b[159:152];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10771_ = b[167:160];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10771_ = b[175:168];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10771_ = b[183:176];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10771_ = b[191:184];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10771_ = b[199:192];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10771_ = b[207:200];
      123'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10771_ = b[215:208];
      123'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10771_ = b[223:216];
      123'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10771_ = b[231:224];
      123'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10771_ = b[239:232];
      123'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10771_ = b[247:240];
      123'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10771_ = b[255:248];
      123'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10771_ = b[263:256];
      123'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10771_ = b[271:264];
      123'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10771_ = b[279:272];
      123'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10771_ = b[287:280];
      123'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10771_ = b[295:288];
      123'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10771_ = b[303:296];
      123'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10771_ = b[311:304];
      123'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10771_ = b[319:312];
      123'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10771_ = b[327:320];
      123'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10771_ = b[335:328];
      123'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10771_ = b[343:336];
      123'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10771_ = b[351:344];
      123'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10771_ = b[359:352];
      123'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10771_ = b[367:360];
      123'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10771_ = b[375:368];
      123'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10771_ = b[383:376];
      123'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10771_ = b[391:384];
      123'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10771_ = b[399:392];
      123'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10771_ = b[407:400];
      123'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10771_ = b[415:408];
      123'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10771_ = b[423:416];
      123'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10771_ = b[431:424];
      123'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10771_ = b[439:432];
      123'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10771_ = b[447:440];
      123'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10771_ = b[455:448];
      123'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10771_ = b[463:456];
      123'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10771_ = b[471:464];
      123'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10771_ = b[479:472];
      123'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10771_ = b[487:480];
      123'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10771_ = b[495:488];
      123'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10771_ = b[503:496];
      123'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10771_ = b[511:504];
      123'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10771_ = b[519:512];
      123'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10771_ = b[527:520];
      123'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10771_ = b[535:528];
      123'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10771_ = b[543:536];
      123'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10771_ = b[551:544];
      123'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10771_ = b[559:552];
      123'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10771_ = b[567:560];
      123'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10771_ = b[575:568];
      123'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10771_ = b[583:576];
      123'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10771_ = b[591:584];
      123'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10771_ = b[599:592];
      123'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10771_ = b[607:600];
      123'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[615:608];
      123'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[623:616];
      123'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[631:624];
      123'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[639:632];
      123'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[647:640];
      123'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[655:648];
      123'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[663:656];
      123'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[671:664];
      123'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[679:672];
      123'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[687:680];
      123'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[695:688];
      123'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[703:696];
      123'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[711:704];
      123'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[719:712];
      123'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[727:720];
      123'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[735:728];
      123'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[743:736];
      123'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[751:744];
      123'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[759:752];
      123'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[767:760];
      123'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[775:768];
      123'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[783:776];
      123'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[791:784];
      123'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[799:792];
      123'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[807:800];
      123'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[815:808];
      123'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[823:816];
      123'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[831:824];
      123'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[839:832];
      123'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[847:840];
      123'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[855:848];
      123'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[863:856];
      123'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[871:864];
      123'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[879:872];
      123'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[887:880];
      123'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[895:888];
      123'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[903:896];
      123'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[911:904];
      123'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[919:912];
      123'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[927:920];
      123'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[935:928];
      123'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[943:936];
      123'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[951:944];
      123'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[959:952];
      123'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[967:960];
      123'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[975:968];
      123'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10771_ = b[983:976];
      default:
        _10771_ = a;
    endcase
  endfunction
  assign vec_data_122 = _10771_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968], data_d1[983:976] }, { _01498_, _01497_, _01496_, _01495_, _01494_, _01493_, _01492_, _01491_, _01490_, _01489_, _01488_, _01487_, _01486_, _01485_, _01484_, _01483_, _01482_, _01481_, _01480_, _01479_, _01478_, _01477_, _01476_, _01475_, _01474_, _01473_, _01472_, _01471_, _01470_, _01469_, _01468_, _01467_, _01466_, _01465_, _01464_, _01463_, _01462_, _01461_, _01460_, _01459_, _01458_, _01457_, _01456_, _01455_, _01454_, _01453_, _01452_, _01451_, _01450_, _01449_, _01448_, _01447_, _01446_, _01445_, _01444_, _01443_, _01442_, _01441_, _01440_, _01439_, _01438_, _01437_, _01436_, _01435_, _01434_, _01433_, _01432_, _01431_, _01430_, _01429_, _01428_, _01427_, _01426_, _01425_, _01424_, _01423_, _01422_, _01421_, _01420_, _01419_, _01418_, _01417_, _01416_, _01415_, _01414_, _01413_, _01412_, _01411_, _01410_, _01409_, _01408_, _01407_, _01406_, _01405_, _01404_, _01403_, _01402_, _01401_, _01400_, _01399_, _01398_, _01397_, _01396_, _01395_, _01394_, _01393_, _01392_, _01391_, _01390_, _01389_, _01388_, _01387_, _01386_, _01385_, _01384_, _01383_, _01382_, _01381_, _01380_, _01379_, _01378_, _01377_, _01376_ });
  assign _01376_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1111011;
  assign _01377_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1111010;
  assign _01378_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1111001;
  assign _01379_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1111000;
  assign _01380_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110111;
  assign _01381_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110110;
  assign _01382_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110101;
  assign _01383_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110100;
  assign _01384_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110011;
  assign _01385_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110010;
  assign _01386_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110001;
  assign _01387_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1110000;
  assign _01388_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101111;
  assign _01389_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101110;
  assign _01390_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101101;
  assign _01391_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101100;
  assign _01392_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101011;
  assign _01393_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101010;
  assign _01394_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101001;
  assign _01395_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1101000;
  assign _01396_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100111;
  assign _01397_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100110;
  assign _01398_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100101;
  assign _01399_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100100;
  assign _01400_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100011;
  assign _01401_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100010;
  assign _01402_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100001;
  assign _01403_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1100000;
  assign _01404_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011111;
  assign _01405_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011110;
  assign _01406_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011101;
  assign _01407_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011100;
  assign _01408_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011011;
  assign _01409_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011010;
  assign _01410_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011001;
  assign _01411_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1011000;
  assign _01412_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010111;
  assign _01413_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010110;
  assign _01414_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010101;
  assign _01415_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010100;
  assign _01416_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010011;
  assign _01417_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010010;
  assign _01418_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010001;
  assign _01419_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1010000;
  assign _01420_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001111;
  assign _01421_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001110;
  assign _01422_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001101;
  assign _01423_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001100;
  assign _01424_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001011;
  assign _01425_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001010;
  assign _01426_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001001;
  assign _01427_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1001000;
  assign _01428_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000111;
  assign _01429_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000110;
  assign _01430_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000101;
  assign _01431_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000100;
  assign _01432_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000011;
  assign _01433_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000010;
  assign _01434_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000001;
  assign _01435_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 7'b1000000;
  assign _01436_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111111;
  assign _01437_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111110;
  assign _01438_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111101;
  assign _01439_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111100;
  assign _01440_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111011;
  assign _01441_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111010;
  assign _01442_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111001;
  assign _01443_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b111000;
  assign _01444_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110111;
  assign _01445_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110110;
  assign _01446_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110101;
  assign _01447_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110100;
  assign _01448_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110011;
  assign _01449_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110010;
  assign _01450_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110001;
  assign _01451_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b110000;
  assign _01452_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101111;
  assign _01453_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101110;
  assign _01454_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101101;
  assign _01455_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101100;
  assign _01456_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101011;
  assign _01457_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101010;
  assign _01458_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101001;
  assign _01459_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12410|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b101000;
  assign _01460_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12409|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100111;
  assign _01461_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100110;
  assign _01462_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100101;
  assign _01463_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100100;
  assign _01464_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100011;
  assign _01465_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100010;
  assign _01466_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100001;
  assign _01467_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 6'b100000;
  assign _01468_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11111;
  assign _01469_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11110;
  assign _01470_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11101;
  assign _01471_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11100;
  assign _01472_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11011;
  assign _01473_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11010;
  assign _01474_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11001;
  assign _01475_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b11000;
  assign _01476_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10111;
  assign _01477_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10110;
  assign _01478_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10101;
  assign _01479_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10100;
  assign _01480_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10011;
  assign _01481_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10010;
  assign _01482_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10001;
  assign _01483_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 5'b10000;
  assign _01484_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1111;
  assign _01485_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1110;
  assign _01486_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1101;
  assign _01487_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1100;
  assign _01488_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1011;
  assign _01489_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1010;
  assign _01490_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1001;
  assign _01491_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 4'b1000;
  assign _01492_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 3'b111;
  assign _01493_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 3'b110;
  assign _01494_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 3'b101;
  assign _01495_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 3'b100;
  assign _01496_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 2'b11;
  assign _01497_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 2'b10;
  assign _01498_ = vec_sum_122_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12370" *) 1'b1;
  function [7:0] _10895_;
    input [7:0] a;
    input [975:0] b;
    input [121:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *)
    (* parallel_case *)
    casez (s)
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _10895_ = b[7:0];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _10895_ = b[15:8];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _10895_ = b[23:16];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _10895_ = b[31:24];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _10895_ = b[39:32];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _10895_ = b[47:40];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _10895_ = b[55:48];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _10895_ = b[63:56];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _10895_ = b[71:64];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _10895_ = b[79:72];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _10895_ = b[87:80];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _10895_ = b[95:88];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _10895_ = b[103:96];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _10895_ = b[111:104];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _10895_ = b[119:112];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _10895_ = b[127:120];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _10895_ = b[135:128];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _10895_ = b[143:136];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _10895_ = b[151:144];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _10895_ = b[159:152];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _10895_ = b[167:160];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _10895_ = b[175:168];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _10895_ = b[183:176];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _10895_ = b[191:184];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _10895_ = b[199:192];
      122'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _10895_ = b[207:200];
      122'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _10895_ = b[215:208];
      122'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _10895_ = b[223:216];
      122'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _10895_ = b[231:224];
      122'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _10895_ = b[239:232];
      122'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _10895_ = b[247:240];
      122'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _10895_ = b[255:248];
      122'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _10895_ = b[263:256];
      122'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _10895_ = b[271:264];
      122'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _10895_ = b[279:272];
      122'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _10895_ = b[287:280];
      122'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _10895_ = b[295:288];
      122'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _10895_ = b[303:296];
      122'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _10895_ = b[311:304];
      122'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _10895_ = b[319:312];
      122'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _10895_ = b[327:320];
      122'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _10895_ = b[335:328];
      122'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _10895_ = b[343:336];
      122'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _10895_ = b[351:344];
      122'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _10895_ = b[359:352];
      122'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _10895_ = b[367:360];
      122'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _10895_ = b[375:368];
      122'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _10895_ = b[383:376];
      122'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _10895_ = b[391:384];
      122'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _10895_ = b[399:392];
      122'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _10895_ = b[407:400];
      122'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _10895_ = b[415:408];
      122'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _10895_ = b[423:416];
      122'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _10895_ = b[431:424];
      122'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _10895_ = b[439:432];
      122'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _10895_ = b[447:440];
      122'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _10895_ = b[455:448];
      122'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _10895_ = b[463:456];
      122'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _10895_ = b[471:464];
      122'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _10895_ = b[479:472];
      122'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _10895_ = b[487:480];
      122'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _10895_ = b[495:488];
      122'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _10895_ = b[503:496];
      122'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _10895_ = b[511:504];
      122'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _10895_ = b[519:512];
      122'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _10895_ = b[527:520];
      122'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _10895_ = b[535:528];
      122'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _10895_ = b[543:536];
      122'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _10895_ = b[551:544];
      122'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _10895_ = b[559:552];
      122'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _10895_ = b[567:560];
      122'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _10895_ = b[575:568];
      122'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _10895_ = b[583:576];
      122'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _10895_ = b[591:584];
      122'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _10895_ = b[599:592];
      122'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _10895_ = b[607:600];
      122'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[615:608];
      122'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[623:616];
      122'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[631:624];
      122'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[639:632];
      122'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[647:640];
      122'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[655:648];
      122'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[663:656];
      122'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[671:664];
      122'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[679:672];
      122'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[687:680];
      122'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[695:688];
      122'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[703:696];
      122'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[711:704];
      122'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[719:712];
      122'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[727:720];
      122'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[735:728];
      122'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[743:736];
      122'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[751:744];
      122'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[759:752];
      122'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[767:760];
      122'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[775:768];
      122'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[783:776];
      122'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[791:784];
      122'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[799:792];
      122'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[807:800];
      122'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[815:808];
      122'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[823:816];
      122'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[831:824];
      122'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[839:832];
      122'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[847:840];
      122'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[855:848];
      122'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[863:856];
      122'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[871:864];
      122'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[879:872];
      122'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[887:880];
      122'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[895:888];
      122'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[903:896];
      122'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[911:904];
      122'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[919:912];
      122'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[927:920];
      122'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[935:928];
      122'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[943:936];
      122'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[951:944];
      122'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[959:952];
      122'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[967:960];
      122'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _10895_ = b[975:968];
      default:
        _10895_ = a;
    endcase
  endfunction
  assign vec_data_121 = _10895_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960], data_d1[975:968] }, { _01620_, _01619_, _01618_, _01617_, _01616_, _01615_, _01614_, _01613_, _01612_, _01611_, _01610_, _01609_, _01608_, _01607_, _01606_, _01605_, _01604_, _01603_, _01602_, _01601_, _01600_, _01599_, _01598_, _01597_, _01596_, _01595_, _01594_, _01593_, _01592_, _01591_, _01590_, _01589_, _01588_, _01587_, _01586_, _01585_, _01584_, _01583_, _01582_, _01581_, _01580_, _01579_, _01578_, _01577_, _01576_, _01575_, _01574_, _01573_, _01572_, _01571_, _01570_, _01569_, _01568_, _01567_, _01566_, _01565_, _01564_, _01563_, _01562_, _01561_, _01560_, _01559_, _01558_, _01557_, _01556_, _01555_, _01554_, _01553_, _01552_, _01551_, _01550_, _01549_, _01548_, _01547_, _01546_, _01545_, _01544_, _01543_, _01542_, _01541_, _01540_, _01539_, _01538_, _01537_, _01536_, _01535_, _01534_, _01533_, _01532_, _01531_, _01530_, _01529_, _01528_, _01527_, _01526_, _01525_, _01524_, _01523_, _01522_, _01521_, _01520_, _01519_, _01518_, _01517_, _01516_, _01515_, _01514_, _01513_, _01512_, _01511_, _01510_, _01509_, _01508_, _01507_, _01506_, _01505_, _01504_, _01503_, _01502_, _01501_, _01500_, _01499_ });
  assign _01499_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1111010;
  assign _01500_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1111001;
  assign _01501_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1111000;
  assign _01502_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110111;
  assign _01503_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110110;
  assign _01504_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110101;
  assign _01505_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110100;
  assign _01506_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110011;
  assign _01507_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110010;
  assign _01508_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110001;
  assign _01509_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1110000;
  assign _01510_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101111;
  assign _01511_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101110;
  assign _01512_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101101;
  assign _01513_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101100;
  assign _01514_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101011;
  assign _01515_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101010;
  assign _01516_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101001;
  assign _01517_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1101000;
  assign _01518_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100111;
  assign _01519_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100110;
  assign _01520_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100101;
  assign _01521_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100100;
  assign _01522_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100011;
  assign _01523_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100010;
  assign _01524_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100001;
  assign _01525_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1100000;
  assign _01526_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011111;
  assign _01527_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011110;
  assign _01528_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011101;
  assign _01529_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011100;
  assign _01530_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011011;
  assign _01531_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011010;
  assign _01532_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011001;
  assign _01533_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1011000;
  assign _01534_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010111;
  assign _01535_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010110;
  assign _01536_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010101;
  assign _01537_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010100;
  assign _01538_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010011;
  assign _01539_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010010;
  assign _01540_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010001;
  assign _01541_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1010000;
  assign _01542_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001111;
  assign _01543_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001110;
  assign _01544_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001101;
  assign _01545_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001100;
  assign _01546_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001011;
  assign _01547_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001010;
  assign _01548_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001001;
  assign _01549_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1001000;
  assign _01550_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000111;
  assign _01551_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000110;
  assign _01552_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000101;
  assign _01553_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000100;
  assign _01554_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000011;
  assign _01555_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000010;
  assign _01556_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000001;
  assign _01557_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 7'b1000000;
  assign _01558_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111111;
  assign _01559_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111110;
  assign _01560_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111101;
  assign _01561_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111100;
  assign _01562_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111011;
  assign _01563_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111010;
  assign _01564_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111001;
  assign _01565_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b111000;
  assign _01566_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110111;
  assign _01567_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110110;
  assign _01568_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110101;
  assign _01569_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110100;
  assign _01570_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110011;
  assign _01571_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110010;
  assign _01572_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110001;
  assign _01573_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b110000;
  assign _01574_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101111;
  assign _01575_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101110;
  assign _01576_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101101;
  assign _01577_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101100;
  assign _01578_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101011;
  assign _01579_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101010;
  assign _01580_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101001;
  assign _01581_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b101000;
  assign _01582_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100111;
  assign _01583_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100110;
  assign _01584_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100101;
  assign _01585_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100100;
  assign _01586_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100011;
  assign _01587_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100010;
  assign _01588_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100001;
  assign _01589_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 6'b100000;
  assign _01590_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11111;
  assign _01591_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11110;
  assign _01592_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11101;
  assign _01593_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11100;
  assign _01594_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11011;
  assign _01595_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11010;
  assign _01596_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11001;
  assign _01597_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b11000;
  assign _01598_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10111;
  assign _01599_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10110;
  assign _01600_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10101;
  assign _01601_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10100;
  assign _01602_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10011;
  assign _01603_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10010;
  assign _01604_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10001;
  assign _01605_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 5'b10000;
  assign _01606_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1111;
  assign _01607_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1110;
  assign _01608_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1101;
  assign _01609_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1100;
  assign _01610_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1011;
  assign _01611_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1010;
  assign _01612_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1001;
  assign _01613_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 4'b1000;
  assign _01614_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 3'b111;
  assign _01615_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 3'b110;
  assign _01616_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 3'b101;
  assign _01617_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 3'b100;
  assign _01618_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 2'b11;
  assign _01619_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 2'b10;
  assign _01620_ = vec_sum_121_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12240" *) 1'b1;
  function [7:0] _11018_;
    input [7:0] a;
    input [967:0] b;
    input [120:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *)
    (* parallel_case *)
    casez (s)
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11018_ = b[7:0];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11018_ = b[15:8];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11018_ = b[23:16];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11018_ = b[31:24];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11018_ = b[39:32];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11018_ = b[47:40];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11018_ = b[55:48];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11018_ = b[63:56];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11018_ = b[71:64];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11018_ = b[79:72];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11018_ = b[87:80];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11018_ = b[95:88];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11018_ = b[103:96];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11018_ = b[111:104];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11018_ = b[119:112];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11018_ = b[127:120];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11018_ = b[135:128];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11018_ = b[143:136];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11018_ = b[151:144];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11018_ = b[159:152];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11018_ = b[167:160];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11018_ = b[175:168];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11018_ = b[183:176];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11018_ = b[191:184];
      121'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11018_ = b[199:192];
      121'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11018_ = b[207:200];
      121'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11018_ = b[215:208];
      121'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11018_ = b[223:216];
      121'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11018_ = b[231:224];
      121'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11018_ = b[239:232];
      121'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11018_ = b[247:240];
      121'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11018_ = b[255:248];
      121'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11018_ = b[263:256];
      121'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11018_ = b[271:264];
      121'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11018_ = b[279:272];
      121'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11018_ = b[287:280];
      121'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11018_ = b[295:288];
      121'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11018_ = b[303:296];
      121'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11018_ = b[311:304];
      121'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11018_ = b[319:312];
      121'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11018_ = b[327:320];
      121'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11018_ = b[335:328];
      121'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11018_ = b[343:336];
      121'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11018_ = b[351:344];
      121'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11018_ = b[359:352];
      121'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11018_ = b[367:360];
      121'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11018_ = b[375:368];
      121'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11018_ = b[383:376];
      121'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11018_ = b[391:384];
      121'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11018_ = b[399:392];
      121'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11018_ = b[407:400];
      121'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11018_ = b[415:408];
      121'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11018_ = b[423:416];
      121'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11018_ = b[431:424];
      121'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11018_ = b[439:432];
      121'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11018_ = b[447:440];
      121'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11018_ = b[455:448];
      121'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11018_ = b[463:456];
      121'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11018_ = b[471:464];
      121'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11018_ = b[479:472];
      121'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11018_ = b[487:480];
      121'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11018_ = b[495:488];
      121'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11018_ = b[503:496];
      121'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11018_ = b[511:504];
      121'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11018_ = b[519:512];
      121'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11018_ = b[527:520];
      121'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11018_ = b[535:528];
      121'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11018_ = b[543:536];
      121'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11018_ = b[551:544];
      121'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11018_ = b[559:552];
      121'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11018_ = b[567:560];
      121'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11018_ = b[575:568];
      121'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11018_ = b[583:576];
      121'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11018_ = b[591:584];
      121'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11018_ = b[599:592];
      121'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11018_ = b[607:600];
      121'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[615:608];
      121'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[623:616];
      121'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[631:624];
      121'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[639:632];
      121'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[647:640];
      121'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[655:648];
      121'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[663:656];
      121'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[671:664];
      121'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[679:672];
      121'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[687:680];
      121'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[695:688];
      121'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[703:696];
      121'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[711:704];
      121'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[719:712];
      121'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[727:720];
      121'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[735:728];
      121'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[743:736];
      121'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[751:744];
      121'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[759:752];
      121'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[767:760];
      121'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[775:768];
      121'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[783:776];
      121'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[791:784];
      121'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[799:792];
      121'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[807:800];
      121'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[815:808];
      121'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[823:816];
      121'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[831:824];
      121'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[839:832];
      121'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[847:840];
      121'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[855:848];
      121'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[863:856];
      121'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[871:864];
      121'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[879:872];
      121'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[887:880];
      121'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[895:888];
      121'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[903:896];
      121'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[911:904];
      121'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[919:912];
      121'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[927:920];
      121'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[935:928];
      121'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[943:936];
      121'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[951:944];
      121'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[959:952];
      121'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11018_ = b[967:960];
      default:
        _11018_ = a;
    endcase
  endfunction
  assign vec_data_120 = _11018_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952], data_d1[967:960] }, { _01741_, _01740_, _01739_, _01738_, _01737_, _01736_, _01735_, _01734_, _01733_, _01732_, _01731_, _01730_, _01729_, _01728_, _01727_, _01726_, _01725_, _01724_, _01723_, _01722_, _01721_, _01720_, _01719_, _01718_, _01717_, _01716_, _01715_, _01714_, _01713_, _01712_, _01711_, _01710_, _01709_, _01708_, _01707_, _01706_, _01705_, _01704_, _01703_, _01702_, _01701_, _01700_, _01699_, _01698_, _01697_, _01696_, _01695_, _01694_, _01693_, _01692_, _01691_, _01690_, _01689_, _01688_, _01687_, _01686_, _01685_, _01684_, _01683_, _01682_, _01681_, _01680_, _01679_, _01678_, _01677_, _01676_, _01675_, _01674_, _01673_, _01672_, _01671_, _01670_, _01669_, _01668_, _01667_, _01666_, _01665_, _01664_, _01663_, _01662_, _01661_, _01660_, _01659_, _01658_, _01657_, _01656_, _01655_, _01654_, _01653_, _01652_, _01651_, _01650_, _01649_, _01648_, _01647_, _01646_, _01645_, _01644_, _01643_, _01642_, _01641_, _01640_, _01639_, _01638_, _01637_, _01636_, _01635_, _01634_, _01633_, _01632_, _01631_, _01630_, _01629_, _01628_, _01627_, _01626_, _01625_, _01624_, _01623_, _01622_, _01621_ });
  assign _01621_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1111001;
  assign _01622_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1111000;
  assign _01623_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110111;
  assign _01624_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110110;
  assign _01625_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110101;
  assign _01626_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110100;
  assign _01627_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110011;
  assign _01628_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110010;
  assign _01629_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110001;
  assign _01630_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1110000;
  assign _01631_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101111;
  assign _01632_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101110;
  assign _01633_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101101;
  assign _01634_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101100;
  assign _01635_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101011;
  assign _01636_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101010;
  assign _01637_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101001;
  assign _01638_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1101000;
  assign _01639_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100111;
  assign _01640_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100110;
  assign _01641_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100101;
  assign _01642_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100100;
  assign _01643_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100011;
  assign _01644_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100010;
  assign _01645_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100001;
  assign _01646_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1100000;
  assign _01647_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011111;
  assign _01648_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011110;
  assign _01649_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011101;
  assign _01650_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011100;
  assign _01651_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011011;
  assign _01652_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011010;
  assign _01653_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011001;
  assign _01654_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1011000;
  assign _01655_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010111;
  assign _01656_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010110;
  assign _01657_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010101;
  assign _01658_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010100;
  assign _01659_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010011;
  assign _01660_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010010;
  assign _01661_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010001;
  assign _01662_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1010000;
  assign _01663_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001111;
  assign _01664_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001110;
  assign _01665_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001101;
  assign _01666_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001100;
  assign _01667_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001011;
  assign _01668_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001010;
  assign _01669_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001001;
  assign _01670_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1001000;
  assign _01671_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000111;
  assign _01672_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000110;
  assign _01673_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000101;
  assign _01674_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000100;
  assign _01675_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000011;
  assign _01676_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000010;
  assign _01677_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12176|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000001;
  assign _01678_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 7'b1000000;
  assign _01679_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111111;
  assign _01680_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111110;
  assign _01681_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111101;
  assign _01682_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111100;
  assign _01683_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111011;
  assign _01684_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111010;
  assign _01685_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111001;
  assign _01686_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b111000;
  assign _01687_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110111;
  assign _01688_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110110;
  assign _01689_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110101;
  assign _01690_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110100;
  assign _01691_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110011;
  assign _01692_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110010;
  assign _01693_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110001;
  assign _01694_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b110000;
  assign _01695_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101111;
  assign _01696_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101110;
  assign _01697_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101101;
  assign _01698_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101100;
  assign _01699_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101011;
  assign _01700_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101010;
  assign _01701_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101001;
  assign _01702_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b101000;
  assign _01703_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100111;
  assign _01704_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100110;
  assign _01705_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100101;
  assign _01706_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100100;
  assign _01707_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100011;
  assign _01708_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100010;
  assign _01709_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100001;
  assign _01710_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 6'b100000;
  assign _01711_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11111;
  assign _01712_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11110;
  assign _01713_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11101;
  assign _01714_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11100;
  assign _01715_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11011;
  assign _01716_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11010;
  assign _01717_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11001;
  assign _01718_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b11000;
  assign _01719_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10111;
  assign _01720_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10110;
  assign _01721_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10101;
  assign _01722_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10100;
  assign _01723_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10011;
  assign _01724_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10010;
  assign _01725_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10001;
  assign _01726_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 5'b10000;
  assign _01727_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1111;
  assign _01728_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1110;
  assign _01729_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1101;
  assign _01730_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1100;
  assign _01731_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1011;
  assign _01732_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1010;
  assign _01733_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1001;
  assign _01734_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 4'b1000;
  assign _01735_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 3'b111;
  assign _01736_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 3'b110;
  assign _01737_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 3'b101;
  assign _01738_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 3'b100;
  assign _01739_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 2'b11;
  assign _01740_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 2'b10;
  assign _01741_ = vec_sum_120_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12111" *) 1'b1;
  function [7:0] _11140_;
    input [7:0] a;
    input [959:0] b;
    input [119:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *)
    (* parallel_case *)
    casez (s)
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11140_ = b[7:0];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11140_ = b[15:8];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11140_ = b[23:16];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11140_ = b[31:24];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11140_ = b[39:32];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11140_ = b[47:40];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11140_ = b[55:48];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11140_ = b[63:56];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11140_ = b[71:64];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11140_ = b[79:72];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11140_ = b[87:80];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11140_ = b[95:88];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11140_ = b[103:96];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11140_ = b[111:104];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11140_ = b[119:112];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11140_ = b[127:120];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11140_ = b[135:128];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11140_ = b[143:136];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11140_ = b[151:144];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11140_ = b[159:152];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11140_ = b[167:160];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11140_ = b[175:168];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11140_ = b[183:176];
      120'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11140_ = b[191:184];
      120'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11140_ = b[199:192];
      120'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11140_ = b[207:200];
      120'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11140_ = b[215:208];
      120'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11140_ = b[223:216];
      120'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11140_ = b[231:224];
      120'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11140_ = b[239:232];
      120'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11140_ = b[247:240];
      120'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11140_ = b[255:248];
      120'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11140_ = b[263:256];
      120'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11140_ = b[271:264];
      120'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11140_ = b[279:272];
      120'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11140_ = b[287:280];
      120'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11140_ = b[295:288];
      120'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11140_ = b[303:296];
      120'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11140_ = b[311:304];
      120'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11140_ = b[319:312];
      120'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11140_ = b[327:320];
      120'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11140_ = b[335:328];
      120'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11140_ = b[343:336];
      120'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11140_ = b[351:344];
      120'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11140_ = b[359:352];
      120'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11140_ = b[367:360];
      120'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11140_ = b[375:368];
      120'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11140_ = b[383:376];
      120'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11140_ = b[391:384];
      120'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11140_ = b[399:392];
      120'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11140_ = b[407:400];
      120'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11140_ = b[415:408];
      120'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11140_ = b[423:416];
      120'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11140_ = b[431:424];
      120'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11140_ = b[439:432];
      120'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11140_ = b[447:440];
      120'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11140_ = b[455:448];
      120'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11140_ = b[463:456];
      120'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11140_ = b[471:464];
      120'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11140_ = b[479:472];
      120'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11140_ = b[487:480];
      120'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11140_ = b[495:488];
      120'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11140_ = b[503:496];
      120'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11140_ = b[511:504];
      120'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11140_ = b[519:512];
      120'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11140_ = b[527:520];
      120'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11140_ = b[535:528];
      120'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11140_ = b[543:536];
      120'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11140_ = b[551:544];
      120'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11140_ = b[559:552];
      120'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11140_ = b[567:560];
      120'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11140_ = b[575:568];
      120'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11140_ = b[583:576];
      120'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11140_ = b[591:584];
      120'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11140_ = b[599:592];
      120'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11140_ = b[607:600];
      120'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[615:608];
      120'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[623:616];
      120'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[631:624];
      120'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[639:632];
      120'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[647:640];
      120'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[655:648];
      120'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[663:656];
      120'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[671:664];
      120'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[679:672];
      120'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[687:680];
      120'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[695:688];
      120'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[703:696];
      120'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[711:704];
      120'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[719:712];
      120'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[727:720];
      120'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[735:728];
      120'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[743:736];
      120'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[751:744];
      120'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[759:752];
      120'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[767:760];
      120'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[775:768];
      120'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[783:776];
      120'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[791:784];
      120'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[799:792];
      120'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[807:800];
      120'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[815:808];
      120'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[823:816];
      120'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[831:824];
      120'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[839:832];
      120'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[847:840];
      120'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[855:848];
      120'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[863:856];
      120'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[871:864];
      120'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[879:872];
      120'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[887:880];
      120'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[895:888];
      120'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[903:896];
      120'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[911:904];
      120'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[919:912];
      120'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[927:920];
      120'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[935:928];
      120'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[943:936];
      120'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[951:944];
      120'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11140_ = b[959:952];
      default:
        _11140_ = a;
    endcase
  endfunction
  assign vec_data_119 = _11140_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944], data_d1[959:952] }, { _01861_, _01860_, _01859_, _01858_, _01857_, _01856_, _01855_, _01854_, _01853_, _01852_, _01851_, _01850_, _01849_, _01848_, _01847_, _01846_, _01845_, _01844_, _01843_, _01842_, _01841_, _01840_, _01839_, _01838_, _01837_, _01836_, _01835_, _01834_, _01833_, _01832_, _01831_, _01830_, _01829_, _01828_, _01827_, _01826_, _01825_, _01824_, _01823_, _01822_, _01821_, _01820_, _01819_, _01818_, _01817_, _01816_, _01815_, _01814_, _01813_, _01812_, _01811_, _01810_, _01809_, _01808_, _01807_, _01806_, _01805_, _01804_, _01803_, _01802_, _01801_, _01800_, _01799_, _01798_, _01797_, _01796_, _01795_, _01794_, _01793_, _01792_, _01791_, _01790_, _01789_, _01788_, _01787_, _01786_, _01785_, _01784_, _01783_, _01782_, _01781_, _01780_, _01779_, _01778_, _01777_, _01776_, _01775_, _01774_, _01773_, _01772_, _01771_, _01770_, _01769_, _01768_, _01767_, _01766_, _01765_, _01764_, _01763_, _01762_, _01761_, _01760_, _01759_, _01758_, _01757_, _01756_, _01755_, _01754_, _01753_, _01752_, _01751_, _01750_, _01749_, _01748_, _01747_, _01746_, _01745_, _01744_, _01743_, _01742_ });
  assign _01742_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1111000;
  assign _01743_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110111;
  assign _01744_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110110;
  assign _01745_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110101;
  assign _01746_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110100;
  assign _01747_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110011;
  assign _01748_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110010;
  assign _01749_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110001;
  assign _01750_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1110000;
  assign _01751_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101111;
  assign _01752_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101110;
  assign _01753_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101101;
  assign _01754_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101100;
  assign _01755_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101011;
  assign _01756_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101010;
  assign _01757_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101001;
  assign _01758_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1101000;
  assign _01759_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100111;
  assign _01760_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100110;
  assign _01761_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100101;
  assign _01762_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100100;
  assign _01763_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100011;
  assign _01764_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100010;
  assign _01765_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100001;
  assign _01766_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1100000;
  assign _01767_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011111;
  assign _01768_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011110;
  assign _01769_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011101;
  assign _01770_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011100;
  assign _01771_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011011;
  assign _01772_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011010;
  assign _01773_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011001;
  assign _01774_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1011000;
  assign _01775_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010111;
  assign _01776_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010110;
  assign _01777_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010101;
  assign _01778_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010100;
  assign _01779_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010011;
  assign _01780_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010010;
  assign _01781_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010001;
  assign _01782_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1010000;
  assign _01783_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001111;
  assign _01784_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001110;
  assign _01785_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001101;
  assign _01786_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001100;
  assign _01787_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001011;
  assign _01788_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001010;
  assign _01789_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001001;
  assign _01790_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1001000;
  assign _01791_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000111;
  assign _01792_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000110;
  assign _01793_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000101;
  assign _01794_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000100;
  assign _01795_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000011;
  assign _01796_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000010;
  assign _01797_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000001;
  assign _01798_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 7'b1000000;
  assign _01799_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111111;
  assign _01800_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111110;
  assign _01801_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111101;
  assign _01802_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111100;
  assign _01803_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111011;
  assign _01804_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111010;
  assign _01805_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111001;
  assign _01806_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b111000;
  assign _01807_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110111;
  assign _01808_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110110;
  assign _01809_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110101;
  assign _01810_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110100;
  assign _01811_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110011;
  assign _01812_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110010;
  assign _01813_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110001;
  assign _01814_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b110000;
  assign _01815_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101111;
  assign _01816_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101110;
  assign _01817_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101101;
  assign _01818_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101100;
  assign _01819_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101011;
  assign _01820_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101010;
  assign _01821_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101001;
  assign _01822_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b101000;
  assign _01823_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100111;
  assign _01824_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100110;
  assign _01825_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100101;
  assign _01826_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100100;
  assign _01827_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100011;
  assign _01828_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100010;
  assign _01829_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100001;
  assign _01830_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 6'b100000;
  assign _01831_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11111;
  assign _01832_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11110;
  assign _01833_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11101;
  assign _01834_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11100;
  assign _01835_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11011;
  assign _01836_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11010;
  assign _01837_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11001;
  assign _01838_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b11000;
  assign _01839_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10111;
  assign _01840_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10110;
  assign _01841_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10101;
  assign _01842_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10100;
  assign _01843_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10011;
  assign _01844_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10010;
  assign _01845_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:12000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10001;
  assign _01846_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 5'b10000;
  assign _01847_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1111;
  assign _01848_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1110;
  assign _01849_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1101;
  assign _01850_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1100;
  assign _01851_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1011;
  assign _01852_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1010;
  assign _01853_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1001;
  assign _01854_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 4'b1000;
  assign _01855_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 3'b111;
  assign _01856_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 3'b110;
  assign _01857_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 3'b101;
  assign _01858_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 3'b100;
  assign _01859_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 2'b11;
  assign _01860_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 2'b10;
  assign _01861_ = vec_sum_119_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11983" *) 1'b1;
  function [7:0] _11261_;
    input [7:0] a;
    input [951:0] b;
    input [118:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *)
    (* parallel_case *)
    casez (s)
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11261_ = b[7:0];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11261_ = b[15:8];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11261_ = b[23:16];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11261_ = b[31:24];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11261_ = b[39:32];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11261_ = b[47:40];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11261_ = b[55:48];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11261_ = b[63:56];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11261_ = b[71:64];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11261_ = b[79:72];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11261_ = b[87:80];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11261_ = b[95:88];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11261_ = b[103:96];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11261_ = b[111:104];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11261_ = b[119:112];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11261_ = b[127:120];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11261_ = b[135:128];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11261_ = b[143:136];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11261_ = b[151:144];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11261_ = b[159:152];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11261_ = b[167:160];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11261_ = b[175:168];
      119'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11261_ = b[183:176];
      119'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11261_ = b[191:184];
      119'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11261_ = b[199:192];
      119'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11261_ = b[207:200];
      119'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11261_ = b[215:208];
      119'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11261_ = b[223:216];
      119'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11261_ = b[231:224];
      119'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11261_ = b[239:232];
      119'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11261_ = b[247:240];
      119'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11261_ = b[255:248];
      119'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11261_ = b[263:256];
      119'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11261_ = b[271:264];
      119'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11261_ = b[279:272];
      119'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11261_ = b[287:280];
      119'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11261_ = b[295:288];
      119'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11261_ = b[303:296];
      119'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11261_ = b[311:304];
      119'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11261_ = b[319:312];
      119'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11261_ = b[327:320];
      119'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11261_ = b[335:328];
      119'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11261_ = b[343:336];
      119'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11261_ = b[351:344];
      119'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11261_ = b[359:352];
      119'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11261_ = b[367:360];
      119'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11261_ = b[375:368];
      119'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11261_ = b[383:376];
      119'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11261_ = b[391:384];
      119'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11261_ = b[399:392];
      119'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11261_ = b[407:400];
      119'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11261_ = b[415:408];
      119'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11261_ = b[423:416];
      119'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11261_ = b[431:424];
      119'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11261_ = b[439:432];
      119'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11261_ = b[447:440];
      119'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11261_ = b[455:448];
      119'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11261_ = b[463:456];
      119'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11261_ = b[471:464];
      119'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11261_ = b[479:472];
      119'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11261_ = b[487:480];
      119'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11261_ = b[495:488];
      119'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11261_ = b[503:496];
      119'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11261_ = b[511:504];
      119'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11261_ = b[519:512];
      119'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11261_ = b[527:520];
      119'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11261_ = b[535:528];
      119'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11261_ = b[543:536];
      119'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11261_ = b[551:544];
      119'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11261_ = b[559:552];
      119'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11261_ = b[567:560];
      119'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11261_ = b[575:568];
      119'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11261_ = b[583:576];
      119'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11261_ = b[591:584];
      119'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11261_ = b[599:592];
      119'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11261_ = b[607:600];
      119'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[615:608];
      119'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[623:616];
      119'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[631:624];
      119'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[639:632];
      119'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[647:640];
      119'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[655:648];
      119'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[663:656];
      119'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[671:664];
      119'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[679:672];
      119'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[687:680];
      119'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[695:688];
      119'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[703:696];
      119'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[711:704];
      119'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[719:712];
      119'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[727:720];
      119'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[735:728];
      119'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[743:736];
      119'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[751:744];
      119'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[759:752];
      119'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[767:760];
      119'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[775:768];
      119'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[783:776];
      119'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[791:784];
      119'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[799:792];
      119'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[807:800];
      119'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[815:808];
      119'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[823:816];
      119'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[831:824];
      119'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[839:832];
      119'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[847:840];
      119'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[855:848];
      119'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[863:856];
      119'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[871:864];
      119'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[879:872];
      119'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[887:880];
      119'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[895:888];
      119'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[903:896];
      119'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[911:904];
      119'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[919:912];
      119'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[927:920];
      119'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[935:928];
      119'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[943:936];
      119'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11261_ = b[951:944];
      default:
        _11261_ = a;
    endcase
  endfunction
  assign vec_data_118 = _11261_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936], data_d1[951:944] }, { _01980_, _01979_, _01978_, _01977_, _01976_, _01975_, _01974_, _01973_, _01972_, _01971_, _01970_, _01969_, _01968_, _01967_, _01966_, _01965_, _01964_, _01963_, _01962_, _01961_, _01960_, _01959_, _01958_, _01957_, _01956_, _01955_, _01954_, _01953_, _01952_, _01951_, _01950_, _01949_, _01948_, _01947_, _01946_, _01945_, _01944_, _01943_, _01942_, _01941_, _01940_, _01939_, _01938_, _01937_, _01936_, _01935_, _01934_, _01933_, _01932_, _01931_, _01930_, _01929_, _01928_, _01927_, _01926_, _01925_, _01924_, _01923_, _01922_, _01921_, _01920_, _01919_, _01918_, _01917_, _01916_, _01915_, _01914_, _01913_, _01912_, _01911_, _01910_, _01909_, _01908_, _01907_, _01906_, _01905_, _01904_, _01903_, _01902_, _01901_, _01900_, _01899_, _01898_, _01897_, _01896_, _01895_, _01894_, _01893_, _01892_, _01891_, _01890_, _01889_, _01888_, _01887_, _01886_, _01885_, _01884_, _01883_, _01882_, _01881_, _01880_, _01879_, _01878_, _01877_, _01876_, _01875_, _01874_, _01873_, _01872_, _01871_, _01870_, _01869_, _01868_, _01867_, _01866_, _01865_, _01864_, _01863_, _01862_ });
  assign _01862_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110111;
  assign _01863_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110110;
  assign _01864_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110101;
  assign _01865_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110100;
  assign _01866_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110011;
  assign _01867_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110010;
  assign _01868_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110001;
  assign _01869_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1110000;
  assign _01870_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101111;
  assign _01871_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101110;
  assign _01872_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101101;
  assign _01873_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101100;
  assign _01874_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101011;
  assign _01875_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101010;
  assign _01876_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101001;
  assign _01877_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1101000;
  assign _01878_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100111;
  assign _01879_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100110;
  assign _01880_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100101;
  assign _01881_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100100;
  assign _01882_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100011;
  assign _01883_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100010;
  assign _01884_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100001;
  assign _01885_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1100000;
  assign _01886_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011111;
  assign _01887_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011110;
  assign _01888_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011101;
  assign _01889_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011100;
  assign _01890_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011011;
  assign _01891_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011010;
  assign _01892_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011001;
  assign _01893_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1011000;
  assign _01894_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010111;
  assign _01895_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010110;
  assign _01896_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010101;
  assign _01897_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010100;
  assign _01898_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010011;
  assign _01899_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010010;
  assign _01900_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010001;
  assign _01901_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1010000;
  assign _01902_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001111;
  assign _01903_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001110;
  assign _01904_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001101;
  assign _01905_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001100;
  assign _01906_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001011;
  assign _01907_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001010;
  assign _01908_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001001;
  assign _01909_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1001000;
  assign _01910_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000111;
  assign _01911_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000110;
  assign _01912_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000101;
  assign _01913_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000100;
  assign _01914_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000011;
  assign _01915_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000010;
  assign _01916_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000001;
  assign _01917_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 7'b1000000;
  assign _01918_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111111;
  assign _01919_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111110;
  assign _01920_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111101;
  assign _01921_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111100;
  assign _01922_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111011;
  assign _01923_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111010;
  assign _01924_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111001;
  assign _01925_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b111000;
  assign _01926_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110111;
  assign _01927_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110110;
  assign _01928_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110101;
  assign _01929_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110100;
  assign _01930_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110011;
  assign _01931_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110010;
  assign _01932_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110001;
  assign _01933_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b110000;
  assign _01934_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101111;
  assign _01935_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101110;
  assign _01936_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101101;
  assign _01937_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101100;
  assign _01938_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101011;
  assign _01939_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101010;
  assign _01940_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101001;
  assign _01941_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b101000;
  assign _01942_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100111;
  assign _01943_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100110;
  assign _01944_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100101;
  assign _01945_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100100;
  assign _01946_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100011;
  assign _01947_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100010;
  assign _01948_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100001;
  assign _01949_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 6'b100000;
  assign _01950_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11111;
  assign _01951_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11110;
  assign _01952_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11101;
  assign _01953_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11100;
  assign _01954_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11011;
  assign _01955_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11010;
  assign _01956_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11001;
  assign _01957_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b11000;
  assign _01958_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10111;
  assign _01959_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10110;
  assign _01960_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10101;
  assign _01961_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10100;
  assign _01962_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10011;
  assign _01963_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10010;
  assign _01964_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10001;
  assign _01965_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 5'b10000;
  assign _01966_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1111;
  assign _01967_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1110;
  assign _01968_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1101;
  assign _01969_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1100;
  assign _01970_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1011;
  assign _01971_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1010;
  assign _01972_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1001;
  assign _01973_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 4'b1000;
  assign _01974_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 3'b111;
  assign _01975_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 3'b110;
  assign _01976_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 3'b101;
  assign _01977_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 3'b100;
  assign _01978_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 2'b11;
  assign _01979_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 2'b10;
  assign _01980_ = vec_sum_118_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11856" *) 1'b1;
  function [7:0] _11381_;
    input [7:0] a;
    input [943:0] b;
    input [117:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *)
    (* parallel_case *)
    casez (s)
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11381_ = b[7:0];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11381_ = b[15:8];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11381_ = b[23:16];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11381_ = b[31:24];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11381_ = b[39:32];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11381_ = b[47:40];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11381_ = b[55:48];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11381_ = b[63:56];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11381_ = b[71:64];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11381_ = b[79:72];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11381_ = b[87:80];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11381_ = b[95:88];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11381_ = b[103:96];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11381_ = b[111:104];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11381_ = b[119:112];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11381_ = b[127:120];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11381_ = b[135:128];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11381_ = b[143:136];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11381_ = b[151:144];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11381_ = b[159:152];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11381_ = b[167:160];
      118'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11381_ = b[175:168];
      118'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11381_ = b[183:176];
      118'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11381_ = b[191:184];
      118'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11381_ = b[199:192];
      118'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11381_ = b[207:200];
      118'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11381_ = b[215:208];
      118'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11381_ = b[223:216];
      118'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11381_ = b[231:224];
      118'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11381_ = b[239:232];
      118'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11381_ = b[247:240];
      118'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11381_ = b[255:248];
      118'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11381_ = b[263:256];
      118'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11381_ = b[271:264];
      118'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11381_ = b[279:272];
      118'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11381_ = b[287:280];
      118'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11381_ = b[295:288];
      118'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11381_ = b[303:296];
      118'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11381_ = b[311:304];
      118'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11381_ = b[319:312];
      118'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11381_ = b[327:320];
      118'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11381_ = b[335:328];
      118'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11381_ = b[343:336];
      118'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11381_ = b[351:344];
      118'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11381_ = b[359:352];
      118'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11381_ = b[367:360];
      118'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11381_ = b[375:368];
      118'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11381_ = b[383:376];
      118'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11381_ = b[391:384];
      118'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11381_ = b[399:392];
      118'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11381_ = b[407:400];
      118'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11381_ = b[415:408];
      118'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11381_ = b[423:416];
      118'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11381_ = b[431:424];
      118'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11381_ = b[439:432];
      118'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11381_ = b[447:440];
      118'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11381_ = b[455:448];
      118'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11381_ = b[463:456];
      118'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11381_ = b[471:464];
      118'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11381_ = b[479:472];
      118'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11381_ = b[487:480];
      118'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11381_ = b[495:488];
      118'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11381_ = b[503:496];
      118'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11381_ = b[511:504];
      118'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11381_ = b[519:512];
      118'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11381_ = b[527:520];
      118'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11381_ = b[535:528];
      118'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11381_ = b[543:536];
      118'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11381_ = b[551:544];
      118'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11381_ = b[559:552];
      118'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11381_ = b[567:560];
      118'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11381_ = b[575:568];
      118'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11381_ = b[583:576];
      118'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11381_ = b[591:584];
      118'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11381_ = b[599:592];
      118'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11381_ = b[607:600];
      118'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[615:608];
      118'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[623:616];
      118'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[631:624];
      118'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[639:632];
      118'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[647:640];
      118'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[655:648];
      118'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[663:656];
      118'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[671:664];
      118'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[679:672];
      118'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[687:680];
      118'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[695:688];
      118'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[703:696];
      118'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[711:704];
      118'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[719:712];
      118'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[727:720];
      118'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[735:728];
      118'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[743:736];
      118'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[751:744];
      118'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[759:752];
      118'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[767:760];
      118'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[775:768];
      118'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[783:776];
      118'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[791:784];
      118'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[799:792];
      118'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[807:800];
      118'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[815:808];
      118'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[823:816];
      118'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[831:824];
      118'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[839:832];
      118'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[847:840];
      118'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[855:848];
      118'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[863:856];
      118'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[871:864];
      118'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[879:872];
      118'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[887:880];
      118'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[895:888];
      118'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[903:896];
      118'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[911:904];
      118'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[919:912];
      118'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[927:920];
      118'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[935:928];
      118'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11381_ = b[943:936];
      default:
        _11381_ = a;
    endcase
  endfunction
  assign vec_data_117 = _11381_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928], data_d1[943:936] }, { _02098_, _02097_, _02096_, _02095_, _02094_, _02093_, _02092_, _02091_, _02090_, _02089_, _02088_, _02087_, _02086_, _02085_, _02084_, _02083_, _02082_, _02081_, _02080_, _02079_, _02078_, _02077_, _02076_, _02075_, _02074_, _02073_, _02072_, _02071_, _02070_, _02069_, _02068_, _02067_, _02066_, _02065_, _02064_, _02063_, _02062_, _02061_, _02060_, _02059_, _02058_, _02057_, _02056_, _02055_, _02054_, _02053_, _02052_, _02051_, _02050_, _02049_, _02048_, _02047_, _02046_, _02045_, _02044_, _02043_, _02042_, _02041_, _02040_, _02039_, _02038_, _02037_, _02036_, _02035_, _02034_, _02033_, _02032_, _02031_, _02030_, _02029_, _02028_, _02027_, _02026_, _02025_, _02024_, _02023_, _02022_, _02021_, _02020_, _02019_, _02018_, _02017_, _02016_, _02015_, _02014_, _02013_, _02012_, _02011_, _02010_, _02009_, _02008_, _02007_, _02006_, _02005_, _02004_, _02003_, _02002_, _02001_, _02000_, _01999_, _01998_, _01997_, _01996_, _01995_, _01994_, _01993_, _01992_, _01991_, _01990_, _01989_, _01988_, _01987_, _01986_, _01985_, _01984_, _01983_, _01982_, _01981_ });
  assign _01981_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110110;
  assign _01982_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110101;
  assign _01983_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110100;
  assign _01984_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110011;
  assign _01985_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110010;
  assign _01986_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110001;
  assign _01987_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1110000;
  assign _01988_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101111;
  assign _01989_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101110;
  assign _01990_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101101;
  assign _01991_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101100;
  assign _01992_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101011;
  assign _01993_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101010;
  assign _01994_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101001;
  assign _01995_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1101000;
  assign _01996_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100111;
  assign _01997_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100110;
  assign _01998_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100101;
  assign _01999_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100100;
  assign _02000_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100011;
  assign _02001_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100010;
  assign _02002_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100001;
  assign _02003_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1100000;
  assign _02004_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011111;
  assign _02005_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011110;
  assign _02006_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011101;
  assign _02007_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011100;
  assign _02008_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011011;
  assign _02009_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011010;
  assign _02010_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011001;
  assign _02011_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1011000;
  assign _02012_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010111;
  assign _02013_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010110;
  assign _02014_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010101;
  assign _02015_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010100;
  assign _02016_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010011;
  assign _02017_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010010;
  assign _02018_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010001;
  assign _02019_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1010000;
  assign _02020_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001111;
  assign _02021_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001110;
  assign _02022_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001101;
  assign _02023_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001100;
  assign _02024_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001011;
  assign _02025_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001010;
  assign _02026_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001001;
  assign _02027_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1001000;
  assign _02028_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000111;
  assign _02029_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000110;
  assign _02030_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000101;
  assign _02031_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000100;
  assign _02032_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000011;
  assign _02033_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000010;
  assign _02034_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000001;
  assign _02035_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 7'b1000000;
  assign _02036_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111111;
  assign _02037_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111110;
  assign _02038_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111101;
  assign _02039_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111100;
  assign _02040_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111011;
  assign _02041_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111010;
  assign _02042_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111001;
  assign _02043_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b111000;
  assign _02044_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110111;
  assign _02045_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110110;
  assign _02046_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110101;
  assign _02047_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110100;
  assign _02048_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110011;
  assign _02049_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110010;
  assign _02050_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110001;
  assign _02051_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b110000;
  assign _02052_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101111;
  assign _02053_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101110;
  assign _02054_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101101;
  assign _02055_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101100;
  assign _02056_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101011;
  assign _02057_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101010;
  assign _02058_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101001;
  assign _02059_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b101000;
  assign _02060_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100111;
  assign _02061_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100110;
  assign _02062_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100101;
  assign _02063_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100100;
  assign _02064_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100011;
  assign _02065_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100010;
  assign _02066_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100001;
  assign _02067_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 6'b100000;
  assign _02068_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11111;
  assign _02069_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11110;
  assign _02070_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11101;
  assign _02071_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11100;
  assign _02072_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11011;
  assign _02073_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11010;
  assign _02074_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11001;
  assign _02075_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b11000;
  assign _02076_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10111;
  assign _02077_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10110;
  assign _02078_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10101;
  assign _02079_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10100;
  assign _02080_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10011;
  assign _02081_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10010;
  assign _02082_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10001;
  assign _02083_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 5'b10000;
  assign _02084_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1111;
  assign _02085_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1110;
  assign _02086_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1101;
  assign _02087_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1100;
  assign _02088_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1011;
  assign _02089_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1010;
  assign _02090_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1001;
  assign _02091_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 4'b1000;
  assign _02092_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 3'b111;
  assign _02093_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 3'b110;
  assign _02094_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 3'b101;
  assign _02095_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 3'b100;
  assign _02096_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 2'b11;
  assign _02097_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 2'b10;
  assign _02098_ = vec_sum_117_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11730" *) 1'b1;
  function [7:0] _11500_;
    input [7:0] a;
    input [935:0] b;
    input [116:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *)
    (* parallel_case *)
    casez (s)
      117'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11500_ = b[7:0];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11500_ = b[15:8];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11500_ = b[23:16];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11500_ = b[31:24];
      117'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11500_ = b[39:32];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11500_ = b[47:40];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11500_ = b[55:48];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11500_ = b[63:56];
      117'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11500_ = b[71:64];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11500_ = b[79:72];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11500_ = b[87:80];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11500_ = b[95:88];
      117'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11500_ = b[103:96];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11500_ = b[111:104];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11500_ = b[119:112];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11500_ = b[127:120];
      117'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11500_ = b[135:128];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11500_ = b[143:136];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11500_ = b[151:144];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11500_ = b[159:152];
      117'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11500_ = b[167:160];
      117'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11500_ = b[175:168];
      117'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11500_ = b[183:176];
      117'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11500_ = b[191:184];
      117'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11500_ = b[199:192];
      117'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11500_ = b[207:200];
      117'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11500_ = b[215:208];
      117'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11500_ = b[223:216];
      117'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11500_ = b[231:224];
      117'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11500_ = b[239:232];
      117'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11500_ = b[247:240];
      117'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11500_ = b[255:248];
      117'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11500_ = b[263:256];
      117'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11500_ = b[271:264];
      117'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11500_ = b[279:272];
      117'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11500_ = b[287:280];
      117'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11500_ = b[295:288];
      117'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11500_ = b[303:296];
      117'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11500_ = b[311:304];
      117'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11500_ = b[319:312];
      117'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11500_ = b[327:320];
      117'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11500_ = b[335:328];
      117'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11500_ = b[343:336];
      117'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11500_ = b[351:344];
      117'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11500_ = b[359:352];
      117'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11500_ = b[367:360];
      117'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11500_ = b[375:368];
      117'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11500_ = b[383:376];
      117'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11500_ = b[391:384];
      117'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11500_ = b[399:392];
      117'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11500_ = b[407:400];
      117'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11500_ = b[415:408];
      117'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11500_ = b[423:416];
      117'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11500_ = b[431:424];
      117'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11500_ = b[439:432];
      117'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11500_ = b[447:440];
      117'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11500_ = b[455:448];
      117'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11500_ = b[463:456];
      117'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11500_ = b[471:464];
      117'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11500_ = b[479:472];
      117'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11500_ = b[487:480];
      117'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11500_ = b[495:488];
      117'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11500_ = b[503:496];
      117'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11500_ = b[511:504];
      117'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11500_ = b[519:512];
      117'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11500_ = b[527:520];
      117'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11500_ = b[535:528];
      117'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11500_ = b[543:536];
      117'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11500_ = b[551:544];
      117'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11500_ = b[559:552];
      117'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11500_ = b[567:560];
      117'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11500_ = b[575:568];
      117'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11500_ = b[583:576];
      117'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11500_ = b[591:584];
      117'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11500_ = b[599:592];
      117'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11500_ = b[607:600];
      117'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[615:608];
      117'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[623:616];
      117'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[631:624];
      117'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[639:632];
      117'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[647:640];
      117'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[655:648];
      117'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[663:656];
      117'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[671:664];
      117'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[679:672];
      117'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[687:680];
      117'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[695:688];
      117'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[703:696];
      117'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[711:704];
      117'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[719:712];
      117'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[727:720];
      117'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[735:728];
      117'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[743:736];
      117'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[751:744];
      117'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[759:752];
      117'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[767:760];
      117'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[775:768];
      117'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[783:776];
      117'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[791:784];
      117'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[799:792];
      117'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[807:800];
      117'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[815:808];
      117'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[823:816];
      117'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[831:824];
      117'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[839:832];
      117'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[847:840];
      117'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[855:848];
      117'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[863:856];
      117'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[871:864];
      117'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[879:872];
      117'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[887:880];
      117'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[895:888];
      117'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[903:896];
      117'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[911:904];
      117'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[919:912];
      117'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[927:920];
      117'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11500_ = b[935:928];
      default:
        _11500_ = a;
    endcase
  endfunction
  assign vec_data_116 = _11500_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920], data_d1[935:928] }, { _02215_, _02214_, _02213_, _02212_, _02211_, _02210_, _02209_, _02208_, _02207_, _02206_, _02205_, _02204_, _02203_, _02202_, _02201_, _02200_, _02199_, _02198_, _02197_, _02196_, _02195_, _02194_, _02193_, _02192_, _02191_, _02190_, _02189_, _02188_, _02187_, _02186_, _02185_, _02184_, _02183_, _02182_, _02181_, _02180_, _02179_, _02178_, _02177_, _02176_, _02175_, _02174_, _02173_, _02172_, _02171_, _02170_, _02169_, _02168_, _02167_, _02166_, _02165_, _02164_, _02163_, _02162_, _02161_, _02160_, _02159_, _02158_, _02157_, _02156_, _02155_, _02154_, _02153_, _02152_, _02151_, _02150_, _02149_, _02148_, _02147_, _02146_, _02145_, _02144_, _02143_, _02142_, _02141_, _02140_, _02139_, _02138_, _02137_, _02136_, _02135_, _02134_, _02133_, _02132_, _02131_, _02130_, _02129_, _02128_, _02127_, _02126_, _02125_, _02124_, _02123_, _02122_, _02121_, _02120_, _02119_, _02118_, _02117_, _02116_, _02115_, _02114_, _02113_, _02112_, _02111_, _02110_, _02109_, _02108_, _02107_, _02106_, _02105_, _02104_, _02103_, _02102_, _02101_, _02100_, _02099_ });
  assign _02099_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110101;
  assign _02100_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110100;
  assign _02101_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110011;
  assign _02102_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110010;
  assign _02103_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110001;
  assign _02104_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1110000;
  assign _02105_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101111;
  assign _02106_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101110;
  assign _02107_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101101;
  assign _02108_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101100;
  assign _02109_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101011;
  assign _02110_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101010;
  assign _02111_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101001;
  assign _02112_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1101000;
  assign _02113_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100111;
  assign _02114_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100110;
  assign _02115_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100101;
  assign _02116_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100100;
  assign _02117_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100011;
  assign _02118_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100010;
  assign _02119_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100001;
  assign _02120_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1100000;
  assign _02121_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011111;
  assign _02122_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011110;
  assign _02123_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011101;
  assign _02124_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011100;
  assign _02125_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011011;
  assign _02126_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011010;
  assign _02127_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011001;
  assign _02128_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1011000;
  assign _02129_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010111;
  assign _02130_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010110;
  assign _02131_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010101;
  assign _02132_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010100;
  assign _02133_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010011;
  assign _02134_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010010;
  assign _02135_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010001;
  assign _02136_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1010000;
  assign _02137_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001111;
  assign _02138_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001110;
  assign _02139_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001101;
  assign _02140_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001100;
  assign _02141_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001011;
  assign _02142_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001010;
  assign _02143_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001001;
  assign _02144_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1001000;
  assign _02145_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000111;
  assign _02146_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000110;
  assign _02147_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000101;
  assign _02148_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000100;
  assign _02149_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000011;
  assign _02150_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000010;
  assign _02151_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000001;
  assign _02152_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 7'b1000000;
  assign _02153_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111111;
  assign _02154_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111110;
  assign _02155_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111101;
  assign _02156_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111100;
  assign _02157_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111011;
  assign _02158_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111010;
  assign _02159_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111001;
  assign _02160_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b111000;
  assign _02161_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110111;
  assign _02162_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110110;
  assign _02163_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110101;
  assign _02164_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110100;
  assign _02165_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110011;
  assign _02166_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110010;
  assign _02167_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110001;
  assign _02168_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b110000;
  assign _02169_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101111;
  assign _02170_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101110;
  assign _02171_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101101;
  assign _02172_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101100;
  assign _02173_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101011;
  assign _02174_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101010;
  assign _02175_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101001;
  assign _02176_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b101000;
  assign _02177_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100111;
  assign _02178_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100110;
  assign _02179_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100101;
  assign _02180_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100100;
  assign _02181_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100011;
  assign _02182_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100010;
  assign _02183_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100001;
  assign _02184_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 6'b100000;
  assign _02185_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11111;
  assign _02186_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11110;
  assign _02187_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11101;
  assign _02188_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11100;
  assign _02189_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11011;
  assign _02190_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11010;
  assign _02191_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11630|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11001;
  assign _02192_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11629|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b11000;
  assign _02193_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11628|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10111;
  assign _02194_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10110;
  assign _02195_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10101;
  assign _02196_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10100;
  assign _02197_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10011;
  assign _02198_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10010;
  assign _02199_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10001;
  assign _02200_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 5'b10000;
  assign _02201_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1111;
  assign _02202_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1110;
  assign _02203_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1101;
  assign _02204_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1100;
  assign _02205_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1011;
  assign _02206_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1010;
  assign _02207_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1001;
  assign _02208_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 4'b1000;
  assign _02209_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 3'b111;
  assign _02210_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 3'b110;
  assign _02211_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 3'b101;
  assign _02212_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 3'b100;
  assign _02213_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 2'b11;
  assign _02214_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 2'b10;
  assign _02215_ = vec_sum_116_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11605" *) 1'b1;
  function [7:0] _11618_;
    input [7:0] a;
    input [927:0] b;
    input [115:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *)
    (* parallel_case *)
    casez (s)
      116'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11618_ = b[7:0];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11618_ = b[15:8];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11618_ = b[23:16];
      116'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11618_ = b[31:24];
      116'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11618_ = b[39:32];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11618_ = b[47:40];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11618_ = b[55:48];
      116'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11618_ = b[63:56];
      116'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11618_ = b[71:64];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11618_ = b[79:72];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11618_ = b[87:80];
      116'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11618_ = b[95:88];
      116'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11618_ = b[103:96];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11618_ = b[111:104];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11618_ = b[119:112];
      116'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11618_ = b[127:120];
      116'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11618_ = b[135:128];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11618_ = b[143:136];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11618_ = b[151:144];
      116'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11618_ = b[159:152];
      116'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11618_ = b[167:160];
      116'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11618_ = b[175:168];
      116'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11618_ = b[183:176];
      116'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11618_ = b[191:184];
      116'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11618_ = b[199:192];
      116'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11618_ = b[207:200];
      116'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11618_ = b[215:208];
      116'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11618_ = b[223:216];
      116'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11618_ = b[231:224];
      116'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11618_ = b[239:232];
      116'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11618_ = b[247:240];
      116'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11618_ = b[255:248];
      116'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11618_ = b[263:256];
      116'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11618_ = b[271:264];
      116'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11618_ = b[279:272];
      116'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11618_ = b[287:280];
      116'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11618_ = b[295:288];
      116'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11618_ = b[303:296];
      116'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11618_ = b[311:304];
      116'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11618_ = b[319:312];
      116'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11618_ = b[327:320];
      116'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11618_ = b[335:328];
      116'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11618_ = b[343:336];
      116'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11618_ = b[351:344];
      116'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11618_ = b[359:352];
      116'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11618_ = b[367:360];
      116'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11618_ = b[375:368];
      116'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11618_ = b[383:376];
      116'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11618_ = b[391:384];
      116'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11618_ = b[399:392];
      116'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11618_ = b[407:400];
      116'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11618_ = b[415:408];
      116'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11618_ = b[423:416];
      116'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11618_ = b[431:424];
      116'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11618_ = b[439:432];
      116'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11618_ = b[447:440];
      116'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11618_ = b[455:448];
      116'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11618_ = b[463:456];
      116'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11618_ = b[471:464];
      116'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11618_ = b[479:472];
      116'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11618_ = b[487:480];
      116'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11618_ = b[495:488];
      116'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11618_ = b[503:496];
      116'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11618_ = b[511:504];
      116'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11618_ = b[519:512];
      116'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11618_ = b[527:520];
      116'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11618_ = b[535:528];
      116'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11618_ = b[543:536];
      116'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11618_ = b[551:544];
      116'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11618_ = b[559:552];
      116'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11618_ = b[567:560];
      116'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11618_ = b[575:568];
      116'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11618_ = b[583:576];
      116'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11618_ = b[591:584];
      116'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11618_ = b[599:592];
      116'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11618_ = b[607:600];
      116'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[615:608];
      116'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[623:616];
      116'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[631:624];
      116'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[639:632];
      116'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[647:640];
      116'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[655:648];
      116'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[663:656];
      116'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[671:664];
      116'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[679:672];
      116'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[687:680];
      116'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[695:688];
      116'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[703:696];
      116'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[711:704];
      116'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[719:712];
      116'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[727:720];
      116'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[735:728];
      116'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[743:736];
      116'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[751:744];
      116'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[759:752];
      116'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[767:760];
      116'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[775:768];
      116'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[783:776];
      116'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[791:784];
      116'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[799:792];
      116'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[807:800];
      116'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[815:808];
      116'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[823:816];
      116'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[831:824];
      116'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[839:832];
      116'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[847:840];
      116'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[855:848];
      116'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[863:856];
      116'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[871:864];
      116'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[879:872];
      116'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[887:880];
      116'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[895:888];
      116'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[903:896];
      116'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[911:904];
      116'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[919:912];
      116'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11618_ = b[927:920];
      default:
        _11618_ = a;
    endcase
  endfunction
  assign vec_data_115 = _11618_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912], data_d1[927:920] }, { _02331_, _02330_, _02329_, _02328_, _02327_, _02326_, _02325_, _02324_, _02323_, _02322_, _02321_, _02320_, _02319_, _02318_, _02317_, _02316_, _02315_, _02314_, _02313_, _02312_, _02311_, _02310_, _02309_, _02308_, _02307_, _02306_, _02305_, _02304_, _02303_, _02302_, _02301_, _02300_, _02299_, _02298_, _02297_, _02296_, _02295_, _02294_, _02293_, _02292_, _02291_, _02290_, _02289_, _02288_, _02287_, _02286_, _02285_, _02284_, _02283_, _02282_, _02281_, _02280_, _02279_, _02278_, _02277_, _02276_, _02275_, _02274_, _02273_, _02272_, _02271_, _02270_, _02269_, _02268_, _02267_, _02266_, _02265_, _02264_, _02263_, _02262_, _02261_, _02260_, _02259_, _02258_, _02257_, _02256_, _02255_, _02254_, _02253_, _02252_, _02251_, _02250_, _02249_, _02248_, _02247_, _02246_, _02245_, _02244_, _02243_, _02242_, _02241_, _02240_, _02239_, _02238_, _02237_, _02236_, _02235_, _02234_, _02233_, _02232_, _02231_, _02230_, _02229_, _02228_, _02227_, _02226_, _02225_, _02224_, _02223_, _02222_, _02221_, _02220_, _02219_, _02218_, _02217_, _02216_ });
  assign _02216_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1110100;
  assign _02217_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1110011;
  assign _02218_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1110010;
  assign _02219_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1110001;
  assign _02220_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1110000;
  assign _02221_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101111;
  assign _02222_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101110;
  assign _02223_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101101;
  assign _02224_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101100;
  assign _02225_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101011;
  assign _02226_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101010;
  assign _02227_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101001;
  assign _02228_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1101000;
  assign _02229_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100111;
  assign _02230_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100110;
  assign _02231_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100101;
  assign _02232_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100100;
  assign _02233_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100011;
  assign _02234_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100010;
  assign _02235_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100001;
  assign _02236_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1100000;
  assign _02237_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011111;
  assign _02238_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011110;
  assign _02239_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011101;
  assign _02240_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011100;
  assign _02241_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011011;
  assign _02242_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011010;
  assign _02243_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011001;
  assign _02244_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1011000;
  assign _02245_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010111;
  assign _02246_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010110;
  assign _02247_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010101;
  assign _02248_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010100;
  assign _02249_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010011;
  assign _02250_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010010;
  assign _02251_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010001;
  assign _02252_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1010000;
  assign _02253_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001111;
  assign _02254_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001110;
  assign _02255_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001101;
  assign _02256_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001100;
  assign _02257_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001011;
  assign _02258_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001010;
  assign _02259_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001001;
  assign _02260_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1001000;
  assign _02261_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000111;
  assign _02262_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000110;
  assign _02263_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000101;
  assign _02264_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000100;
  assign _02265_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000011;
  assign _02266_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000010;
  assign _02267_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000001;
  assign _02268_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 7'b1000000;
  assign _02269_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111111;
  assign _02270_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111110;
  assign _02271_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111101;
  assign _02272_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111100;
  assign _02273_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111011;
  assign _02274_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111010;
  assign _02275_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111001;
  assign _02276_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b111000;
  assign _02277_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110111;
  assign _02278_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110110;
  assign _02279_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110101;
  assign _02280_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110100;
  assign _02281_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110011;
  assign _02282_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110010;
  assign _02283_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110001;
  assign _02284_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b110000;
  assign _02285_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101111;
  assign _02286_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101110;
  assign _02287_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101101;
  assign _02288_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101100;
  assign _02289_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101011;
  assign _02290_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101010;
  assign _02291_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101001;
  assign _02292_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b101000;
  assign _02293_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100111;
  assign _02294_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100110;
  assign _02295_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100101;
  assign _02296_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100100;
  assign _02297_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100011;
  assign _02298_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100010;
  assign _02299_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100001;
  assign _02300_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 6'b100000;
  assign _02301_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11111;
  assign _02302_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11110;
  assign _02303_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11101;
  assign _02304_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11100;
  assign _02305_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11011;
  assign _02306_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11010;
  assign _02307_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11001;
  assign _02308_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b11000;
  assign _02309_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10111;
  assign _02310_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10110;
  assign _02311_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10101;
  assign _02312_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10100;
  assign _02313_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10011;
  assign _02314_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10010;
  assign _02315_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10001;
  assign _02316_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 5'b10000;
  assign _02317_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1111;
  assign _02318_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1110;
  assign _02319_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1101;
  assign _02320_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1100;
  assign _02321_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1011;
  assign _02322_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1010;
  assign _02323_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1001;
  assign _02324_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 4'b1000;
  assign _02325_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 3'b111;
  assign _02326_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 3'b110;
  assign _02327_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 3'b101;
  assign _02328_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 3'b100;
  assign _02329_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 2'b11;
  assign _02330_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 2'b10;
  assign _02331_ = vec_sum_115_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11481" *) 1'b1;
  function [7:0] _11735_;
    input [7:0] a;
    input [919:0] b;
    input [114:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *)
    (* parallel_case *)
    casez (s)
      115'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11735_ = b[7:0];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11735_ = b[15:8];
      115'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11735_ = b[23:16];
      115'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11735_ = b[31:24];
      115'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11735_ = b[39:32];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11735_ = b[47:40];
      115'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11735_ = b[55:48];
      115'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11735_ = b[63:56];
      115'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11735_ = b[71:64];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11735_ = b[79:72];
      115'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11735_ = b[87:80];
      115'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11735_ = b[95:88];
      115'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11735_ = b[103:96];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11735_ = b[111:104];
      115'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11735_ = b[119:112];
      115'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11735_ = b[127:120];
      115'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11735_ = b[135:128];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11735_ = b[143:136];
      115'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11735_ = b[151:144];
      115'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11735_ = b[159:152];
      115'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11735_ = b[167:160];
      115'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11735_ = b[175:168];
      115'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11735_ = b[183:176];
      115'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11735_ = b[191:184];
      115'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11735_ = b[199:192];
      115'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11735_ = b[207:200];
      115'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11735_ = b[215:208];
      115'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11735_ = b[223:216];
      115'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11735_ = b[231:224];
      115'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11735_ = b[239:232];
      115'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11735_ = b[247:240];
      115'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11735_ = b[255:248];
      115'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11735_ = b[263:256];
      115'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11735_ = b[271:264];
      115'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11735_ = b[279:272];
      115'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11735_ = b[287:280];
      115'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11735_ = b[295:288];
      115'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11735_ = b[303:296];
      115'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11735_ = b[311:304];
      115'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11735_ = b[319:312];
      115'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11735_ = b[327:320];
      115'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11735_ = b[335:328];
      115'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11735_ = b[343:336];
      115'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11735_ = b[351:344];
      115'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11735_ = b[359:352];
      115'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11735_ = b[367:360];
      115'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11735_ = b[375:368];
      115'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11735_ = b[383:376];
      115'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11735_ = b[391:384];
      115'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11735_ = b[399:392];
      115'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11735_ = b[407:400];
      115'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11735_ = b[415:408];
      115'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11735_ = b[423:416];
      115'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11735_ = b[431:424];
      115'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11735_ = b[439:432];
      115'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11735_ = b[447:440];
      115'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11735_ = b[455:448];
      115'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11735_ = b[463:456];
      115'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11735_ = b[471:464];
      115'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11735_ = b[479:472];
      115'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11735_ = b[487:480];
      115'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11735_ = b[495:488];
      115'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11735_ = b[503:496];
      115'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11735_ = b[511:504];
      115'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11735_ = b[519:512];
      115'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11735_ = b[527:520];
      115'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11735_ = b[535:528];
      115'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11735_ = b[543:536];
      115'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11735_ = b[551:544];
      115'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11735_ = b[559:552];
      115'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11735_ = b[567:560];
      115'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11735_ = b[575:568];
      115'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11735_ = b[583:576];
      115'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11735_ = b[591:584];
      115'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11735_ = b[599:592];
      115'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11735_ = b[607:600];
      115'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[615:608];
      115'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[623:616];
      115'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[631:624];
      115'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[639:632];
      115'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[647:640];
      115'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[655:648];
      115'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[663:656];
      115'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[671:664];
      115'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[679:672];
      115'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[687:680];
      115'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[695:688];
      115'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[703:696];
      115'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[711:704];
      115'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[719:712];
      115'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[727:720];
      115'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[735:728];
      115'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[743:736];
      115'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[751:744];
      115'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[759:752];
      115'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[767:760];
      115'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[775:768];
      115'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[783:776];
      115'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[791:784];
      115'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[799:792];
      115'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[807:800];
      115'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[815:808];
      115'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[823:816];
      115'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[831:824];
      115'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[839:832];
      115'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[847:840];
      115'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[855:848];
      115'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[863:856];
      115'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[871:864];
      115'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[879:872];
      115'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[887:880];
      115'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[895:888];
      115'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[903:896];
      115'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[911:904];
      115'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11735_ = b[919:912];
      default:
        _11735_ = a;
    endcase
  endfunction
  assign vec_data_114 = _11735_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904], data_d1[919:912] }, { _02446_, _02445_, _02444_, _02443_, _02442_, _02441_, _02440_, _02439_, _02438_, _02437_, _02436_, _02435_, _02434_, _02433_, _02432_, _02431_, _02430_, _02429_, _02428_, _02427_, _02426_, _02425_, _02424_, _02423_, _02422_, _02421_, _02420_, _02419_, _02418_, _02417_, _02416_, _02415_, _02414_, _02413_, _02412_, _02411_, _02410_, _02409_, _02408_, _02407_, _02406_, _02405_, _02404_, _02403_, _02402_, _02401_, _02400_, _02399_, _02398_, _02397_, _02396_, _02395_, _02394_, _02393_, _02392_, _02391_, _02390_, _02389_, _02388_, _02387_, _02386_, _02385_, _02384_, _02383_, _02382_, _02381_, _02380_, _02379_, _02378_, _02377_, _02376_, _02375_, _02374_, _02373_, _02372_, _02371_, _02370_, _02369_, _02368_, _02367_, _02366_, _02365_, _02364_, _02363_, _02362_, _02361_, _02360_, _02359_, _02358_, _02357_, _02356_, _02355_, _02354_, _02353_, _02352_, _02351_, _02350_, _02349_, _02348_, _02347_, _02346_, _02345_, _02344_, _02343_, _02342_, _02341_, _02340_, _02339_, _02338_, _02337_, _02336_, _02335_, _02334_, _02333_, _02332_ });
  assign _02332_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1110011;
  assign _02333_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1110010;
  assign _02334_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1110001;
  assign _02335_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1110000;
  assign _02336_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101111;
  assign _02337_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101110;
  assign _02338_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101101;
  assign _02339_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101100;
  assign _02340_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101011;
  assign _02341_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101010;
  assign _02342_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101001;
  assign _02343_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1101000;
  assign _02344_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100111;
  assign _02345_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100110;
  assign _02346_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100101;
  assign _02347_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100100;
  assign _02348_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100011;
  assign _02349_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100010;
  assign _02350_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100001;
  assign _02351_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1100000;
  assign _02352_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011111;
  assign _02353_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011110;
  assign _02354_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011101;
  assign _02355_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011100;
  assign _02356_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011011;
  assign _02357_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011010;
  assign _02358_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011001;
  assign _02359_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1011000;
  assign _02360_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010111;
  assign _02361_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010110;
  assign _02362_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010101;
  assign _02363_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010100;
  assign _02364_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010011;
  assign _02365_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010010;
  assign _02366_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010001;
  assign _02367_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1010000;
  assign _02368_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001111;
  assign _02369_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001110;
  assign _02370_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001101;
  assign _02371_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001100;
  assign _02372_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001011;
  assign _02373_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001010;
  assign _02374_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001001;
  assign _02375_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1001000;
  assign _02376_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000111;
  assign _02377_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000110;
  assign _02378_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000101;
  assign _02379_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000100;
  assign _02380_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000011;
  assign _02381_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000010;
  assign _02382_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000001;
  assign _02383_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 7'b1000000;
  assign _02384_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111111;
  assign _02385_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111110;
  assign _02386_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111101;
  assign _02387_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111100;
  assign _02388_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111011;
  assign _02389_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111010;
  assign _02390_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111001;
  assign _02391_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b111000;
  assign _02392_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110111;
  assign _02393_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110110;
  assign _02394_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110101;
  assign _02395_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11410|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110100;
  assign _02396_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11409|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110011;
  assign _02397_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110010;
  assign _02398_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110001;
  assign _02399_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b110000;
  assign _02400_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101111;
  assign _02401_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101110;
  assign _02402_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101101;
  assign _02403_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101100;
  assign _02404_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101011;
  assign _02405_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101010;
  assign _02406_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101001;
  assign _02407_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b101000;
  assign _02408_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100111;
  assign _02409_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100110;
  assign _02410_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100101;
  assign _02411_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100100;
  assign _02412_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100011;
  assign _02413_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100010;
  assign _02414_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100001;
  assign _02415_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 6'b100000;
  assign _02416_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11111;
  assign _02417_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11110;
  assign _02418_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11101;
  assign _02419_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11100;
  assign _02420_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11011;
  assign _02421_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11010;
  assign _02422_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11001;
  assign _02423_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b11000;
  assign _02424_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10111;
  assign _02425_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10110;
  assign _02426_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10101;
  assign _02427_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10100;
  assign _02428_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10011;
  assign _02429_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10010;
  assign _02430_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10001;
  assign _02431_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 5'b10000;
  assign _02432_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1111;
  assign _02433_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1110;
  assign _02434_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1101;
  assign _02435_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1100;
  assign _02436_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1011;
  assign _02437_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1010;
  assign _02438_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1001;
  assign _02439_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 4'b1000;
  assign _02440_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 3'b111;
  assign _02441_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 3'b110;
  assign _02442_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 3'b101;
  assign _02443_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 3'b100;
  assign _02444_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 2'b11;
  assign _02445_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 2'b10;
  assign _02446_ = vec_sum_114_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11358" *) 1'b1;
  function [7:0] _11851_;
    input [7:0] a;
    input [911:0] b;
    input [113:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *)
    (* parallel_case *)
    casez (s)
      114'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11851_ = b[7:0];
      114'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11851_ = b[15:8];
      114'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11851_ = b[23:16];
      114'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11851_ = b[31:24];
      114'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11851_ = b[39:32];
      114'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11851_ = b[47:40];
      114'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11851_ = b[55:48];
      114'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11851_ = b[63:56];
      114'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11851_ = b[71:64];
      114'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11851_ = b[79:72];
      114'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11851_ = b[87:80];
      114'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11851_ = b[95:88];
      114'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11851_ = b[103:96];
      114'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11851_ = b[111:104];
      114'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11851_ = b[119:112];
      114'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11851_ = b[127:120];
      114'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11851_ = b[135:128];
      114'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11851_ = b[143:136];
      114'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11851_ = b[151:144];
      114'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11851_ = b[159:152];
      114'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11851_ = b[167:160];
      114'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11851_ = b[175:168];
      114'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11851_ = b[183:176];
      114'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11851_ = b[191:184];
      114'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11851_ = b[199:192];
      114'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11851_ = b[207:200];
      114'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11851_ = b[215:208];
      114'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11851_ = b[223:216];
      114'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11851_ = b[231:224];
      114'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11851_ = b[239:232];
      114'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11851_ = b[247:240];
      114'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11851_ = b[255:248];
      114'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11851_ = b[263:256];
      114'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11851_ = b[271:264];
      114'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11851_ = b[279:272];
      114'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11851_ = b[287:280];
      114'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11851_ = b[295:288];
      114'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11851_ = b[303:296];
      114'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11851_ = b[311:304];
      114'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11851_ = b[319:312];
      114'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11851_ = b[327:320];
      114'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11851_ = b[335:328];
      114'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11851_ = b[343:336];
      114'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11851_ = b[351:344];
      114'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11851_ = b[359:352];
      114'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11851_ = b[367:360];
      114'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11851_ = b[375:368];
      114'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11851_ = b[383:376];
      114'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11851_ = b[391:384];
      114'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11851_ = b[399:392];
      114'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11851_ = b[407:400];
      114'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11851_ = b[415:408];
      114'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11851_ = b[423:416];
      114'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11851_ = b[431:424];
      114'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11851_ = b[439:432];
      114'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11851_ = b[447:440];
      114'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11851_ = b[455:448];
      114'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11851_ = b[463:456];
      114'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11851_ = b[471:464];
      114'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11851_ = b[479:472];
      114'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11851_ = b[487:480];
      114'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11851_ = b[495:488];
      114'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11851_ = b[503:496];
      114'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11851_ = b[511:504];
      114'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11851_ = b[519:512];
      114'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11851_ = b[527:520];
      114'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11851_ = b[535:528];
      114'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11851_ = b[543:536];
      114'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11851_ = b[551:544];
      114'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11851_ = b[559:552];
      114'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11851_ = b[567:560];
      114'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11851_ = b[575:568];
      114'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11851_ = b[583:576];
      114'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11851_ = b[591:584];
      114'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11851_ = b[599:592];
      114'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11851_ = b[607:600];
      114'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[615:608];
      114'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[623:616];
      114'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[631:624];
      114'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[639:632];
      114'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[647:640];
      114'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[655:648];
      114'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[663:656];
      114'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[671:664];
      114'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[679:672];
      114'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[687:680];
      114'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[695:688];
      114'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[703:696];
      114'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[711:704];
      114'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[719:712];
      114'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[727:720];
      114'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[735:728];
      114'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[743:736];
      114'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[751:744];
      114'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[759:752];
      114'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[767:760];
      114'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[775:768];
      114'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[783:776];
      114'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[791:784];
      114'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[799:792];
      114'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[807:800];
      114'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[815:808];
      114'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[823:816];
      114'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[831:824];
      114'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[839:832];
      114'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[847:840];
      114'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[855:848];
      114'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[863:856];
      114'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[871:864];
      114'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[879:872];
      114'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[887:880];
      114'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[895:888];
      114'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[903:896];
      114'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11851_ = b[911:904];
      default:
        _11851_ = a;
    endcase
  endfunction
  assign vec_data_113 = _11851_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896], data_d1[911:904] }, { _02560_, _02559_, _02558_, _02557_, _02556_, _02555_, _02554_, _02553_, _02552_, _02551_, _02550_, _02549_, _02548_, _02547_, _02546_, _02545_, _02544_, _02543_, _02542_, _02541_, _02540_, _02539_, _02538_, _02537_, _02536_, _02535_, _02534_, _02533_, _02532_, _02531_, _02530_, _02529_, _02528_, _02527_, _02526_, _02525_, _02524_, _02523_, _02522_, _02521_, _02520_, _02519_, _02518_, _02517_, _02516_, _02515_, _02514_, _02513_, _02512_, _02511_, _02510_, _02509_, _02508_, _02507_, _02506_, _02505_, _02504_, _02503_, _02502_, _02501_, _02500_, _02499_, _02498_, _02497_, _02496_, _02495_, _02494_, _02493_, _02492_, _02491_, _02490_, _02489_, _02488_, _02487_, _02486_, _02485_, _02484_, _02483_, _02482_, _02481_, _02480_, _02479_, _02478_, _02477_, _02476_, _02475_, _02474_, _02473_, _02472_, _02471_, _02470_, _02469_, _02468_, _02467_, _02466_, _02465_, _02464_, _02463_, _02462_, _02461_, _02460_, _02459_, _02458_, _02457_, _02456_, _02455_, _02454_, _02453_, _02452_, _02451_, _02450_, _02449_, _02448_, _02447_ });
  assign _02447_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1110010;
  assign _02448_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1110001;
  assign _02449_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1110000;
  assign _02450_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101111;
  assign _02451_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101110;
  assign _02452_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101101;
  assign _02453_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101100;
  assign _02454_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101011;
  assign _02455_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101010;
  assign _02456_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101001;
  assign _02457_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1101000;
  assign _02458_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100111;
  assign _02459_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100110;
  assign _02460_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100101;
  assign _02461_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100100;
  assign _02462_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100011;
  assign _02463_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100010;
  assign _02464_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100001;
  assign _02465_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1100000;
  assign _02466_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011111;
  assign _02467_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011110;
  assign _02468_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011101;
  assign _02469_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011100;
  assign _02470_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011011;
  assign _02471_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011010;
  assign _02472_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011001;
  assign _02473_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1011000;
  assign _02474_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010111;
  assign _02475_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010110;
  assign _02476_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010101;
  assign _02477_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010100;
  assign _02478_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010011;
  assign _02479_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010010;
  assign _02480_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010001;
  assign _02481_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1010000;
  assign _02482_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001111;
  assign _02483_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001110;
  assign _02484_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001101;
  assign _02485_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001100;
  assign _02486_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001011;
  assign _02487_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001010;
  assign _02488_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001001;
  assign _02489_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1001000;
  assign _02490_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000111;
  assign _02491_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000110;
  assign _02492_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000101;
  assign _02493_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000100;
  assign _02494_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000011;
  assign _02495_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000010;
  assign _02496_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000001;
  assign _02497_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 7'b1000000;
  assign _02498_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111111;
  assign _02499_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111110;
  assign _02500_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111101;
  assign _02501_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111100;
  assign _02502_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111011;
  assign _02503_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111010;
  assign _02504_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111001;
  assign _02505_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b111000;
  assign _02506_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110111;
  assign _02507_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110110;
  assign _02508_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110101;
  assign _02509_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110100;
  assign _02510_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110011;
  assign _02511_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110010;
  assign _02512_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110001;
  assign _02513_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b110000;
  assign _02514_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101111;
  assign _02515_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101110;
  assign _02516_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101101;
  assign _02517_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101100;
  assign _02518_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101011;
  assign _02519_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101010;
  assign _02520_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101001;
  assign _02521_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b101000;
  assign _02522_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100111;
  assign _02523_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100110;
  assign _02524_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100101;
  assign _02525_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100100;
  assign _02526_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100011;
  assign _02527_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100010;
  assign _02528_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100001;
  assign _02529_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 6'b100000;
  assign _02530_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11111;
  assign _02531_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11110;
  assign _02532_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11101;
  assign _02533_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11100;
  assign _02534_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11011;
  assign _02535_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11010;
  assign _02536_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11001;
  assign _02537_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b11000;
  assign _02538_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10111;
  assign _02539_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10110;
  assign _02540_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10101;
  assign _02541_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10100;
  assign _02542_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10011;
  assign _02543_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10010;
  assign _02544_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10001;
  assign _02545_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 5'b10000;
  assign _02546_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1111;
  assign _02547_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1110;
  assign _02548_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1101;
  assign _02549_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1100;
  assign _02550_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1011;
  assign _02551_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1010;
  assign _02552_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1001;
  assign _02553_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 4'b1000;
  assign _02554_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 3'b111;
  assign _02555_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 3'b110;
  assign _02556_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 3'b101;
  assign _02557_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 3'b100;
  assign _02558_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 2'b11;
  assign _02559_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 2'b10;
  assign _02560_ = vec_sum_113_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11236" *) 1'b1;
  function [7:0] _11966_;
    input [7:0] a;
    input [903:0] b;
    input [112:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *)
    (* parallel_case *)
    casez (s)
      113'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _11966_ = b[7:0];
      113'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _11966_ = b[15:8];
      113'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _11966_ = b[23:16];
      113'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _11966_ = b[31:24];
      113'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _11966_ = b[39:32];
      113'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _11966_ = b[47:40];
      113'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _11966_ = b[55:48];
      113'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _11966_ = b[63:56];
      113'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _11966_ = b[71:64];
      113'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _11966_ = b[79:72];
      113'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _11966_ = b[87:80];
      113'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _11966_ = b[95:88];
      113'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _11966_ = b[103:96];
      113'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _11966_ = b[111:104];
      113'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _11966_ = b[119:112];
      113'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _11966_ = b[127:120];
      113'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _11966_ = b[135:128];
      113'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _11966_ = b[143:136];
      113'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _11966_ = b[151:144];
      113'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _11966_ = b[159:152];
      113'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _11966_ = b[167:160];
      113'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _11966_ = b[175:168];
      113'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _11966_ = b[183:176];
      113'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _11966_ = b[191:184];
      113'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _11966_ = b[199:192];
      113'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _11966_ = b[207:200];
      113'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _11966_ = b[215:208];
      113'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _11966_ = b[223:216];
      113'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _11966_ = b[231:224];
      113'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _11966_ = b[239:232];
      113'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _11966_ = b[247:240];
      113'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _11966_ = b[255:248];
      113'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _11966_ = b[263:256];
      113'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _11966_ = b[271:264];
      113'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _11966_ = b[279:272];
      113'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _11966_ = b[287:280];
      113'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _11966_ = b[295:288];
      113'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _11966_ = b[303:296];
      113'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _11966_ = b[311:304];
      113'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _11966_ = b[319:312];
      113'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _11966_ = b[327:320];
      113'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _11966_ = b[335:328];
      113'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _11966_ = b[343:336];
      113'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _11966_ = b[351:344];
      113'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _11966_ = b[359:352];
      113'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _11966_ = b[367:360];
      113'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _11966_ = b[375:368];
      113'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _11966_ = b[383:376];
      113'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _11966_ = b[391:384];
      113'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _11966_ = b[399:392];
      113'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _11966_ = b[407:400];
      113'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _11966_ = b[415:408];
      113'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _11966_ = b[423:416];
      113'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _11966_ = b[431:424];
      113'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _11966_ = b[439:432];
      113'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _11966_ = b[447:440];
      113'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _11966_ = b[455:448];
      113'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _11966_ = b[463:456];
      113'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _11966_ = b[471:464];
      113'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _11966_ = b[479:472];
      113'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _11966_ = b[487:480];
      113'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _11966_ = b[495:488];
      113'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _11966_ = b[503:496];
      113'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _11966_ = b[511:504];
      113'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _11966_ = b[519:512];
      113'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _11966_ = b[527:520];
      113'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _11966_ = b[535:528];
      113'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _11966_ = b[543:536];
      113'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _11966_ = b[551:544];
      113'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _11966_ = b[559:552];
      113'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _11966_ = b[567:560];
      113'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _11966_ = b[575:568];
      113'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _11966_ = b[583:576];
      113'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _11966_ = b[591:584];
      113'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _11966_ = b[599:592];
      113'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _11966_ = b[607:600];
      113'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[615:608];
      113'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[623:616];
      113'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[631:624];
      113'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[639:632];
      113'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[647:640];
      113'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[655:648];
      113'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[663:656];
      113'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[671:664];
      113'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[679:672];
      113'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[687:680];
      113'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[695:688];
      113'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[703:696];
      113'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[711:704];
      113'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[719:712];
      113'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[727:720];
      113'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[735:728];
      113'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[743:736];
      113'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[751:744];
      113'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[759:752];
      113'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[767:760];
      113'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[775:768];
      113'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[783:776];
      113'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[791:784];
      113'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[799:792];
      113'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[807:800];
      113'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[815:808];
      113'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[823:816];
      113'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[831:824];
      113'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[839:832];
      113'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[847:840];
      113'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[855:848];
      113'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[863:856];
      113'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[871:864];
      113'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[879:872];
      113'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[887:880];
      113'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[895:888];
      113'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _11966_ = b[903:896];
      default:
        _11966_ = a;
    endcase
  endfunction
  assign vec_data_112 = _11966_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888], data_d1[903:896] }, { _02673_, _02672_, _02671_, _02670_, _02669_, _02668_, _02667_, _02666_, _02665_, _02664_, _02663_, _02662_, _02661_, _02660_, _02659_, _02658_, _02657_, _02656_, _02655_, _02654_, _02653_, _02652_, _02651_, _02650_, _02649_, _02648_, _02647_, _02646_, _02645_, _02644_, _02643_, _02642_, _02641_, _02640_, _02639_, _02638_, _02637_, _02636_, _02635_, _02634_, _02633_, _02632_, _02631_, _02630_, _02629_, _02628_, _02627_, _02626_, _02625_, _02624_, _02623_, _02622_, _02621_, _02620_, _02619_, _02618_, _02617_, _02616_, _02615_, _02614_, _02613_, _02612_, _02611_, _02610_, _02609_, _02608_, _02607_, _02606_, _02605_, _02604_, _02603_, _02602_, _02601_, _02600_, _02599_, _02598_, _02597_, _02596_, _02595_, _02594_, _02593_, _02592_, _02591_, _02590_, _02589_, _02588_, _02587_, _02586_, _02585_, _02584_, _02583_, _02582_, _02581_, _02580_, _02579_, _02578_, _02577_, _02576_, _02575_, _02574_, _02573_, _02572_, _02571_, _02570_, _02569_, _02568_, _02567_, _02566_, _02565_, _02564_, _02563_, _02562_, _02561_ });
  assign _02561_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1110001;
  assign _02562_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1110000;
  assign _02563_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101111;
  assign _02564_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101110;
  assign _02565_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101101;
  assign _02566_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101100;
  assign _02567_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101011;
  assign _02568_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101010;
  assign _02569_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101001;
  assign _02570_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1101000;
  assign _02571_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100111;
  assign _02572_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100110;
  assign _02573_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100101;
  assign _02574_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100100;
  assign _02575_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100011;
  assign _02576_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100010;
  assign _02577_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100001;
  assign _02578_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1100000;
  assign _02579_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011111;
  assign _02580_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011110;
  assign _02581_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011101;
  assign _02582_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011100;
  assign _02583_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011011;
  assign _02584_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011010;
  assign _02585_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011001;
  assign _02586_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1011000;
  assign _02587_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010111;
  assign _02588_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010110;
  assign _02589_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010101;
  assign _02590_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010100;
  assign _02591_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010011;
  assign _02592_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010010;
  assign _02593_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010001;
  assign _02594_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1010000;
  assign _02595_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001111;
  assign _02596_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001110;
  assign _02597_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001101;
  assign _02598_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001100;
  assign _02599_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001011;
  assign _02600_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001010;
  assign _02601_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001001;
  assign _02602_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1001000;
  assign _02603_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000111;
  assign _02604_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000110;
  assign _02605_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000101;
  assign _02606_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000100;
  assign _02607_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000011;
  assign _02608_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000010;
  assign _02609_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000001;
  assign _02610_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 7'b1000000;
  assign _02611_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111111;
  assign _02612_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111110;
  assign _02613_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11176|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111101;
  assign _02614_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111100;
  assign _02615_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111011;
  assign _02616_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111010;
  assign _02617_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111001;
  assign _02618_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b111000;
  assign _02619_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110111;
  assign _02620_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110110;
  assign _02621_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110101;
  assign _02622_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110100;
  assign _02623_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110011;
  assign _02624_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110010;
  assign _02625_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110001;
  assign _02626_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b110000;
  assign _02627_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101111;
  assign _02628_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101110;
  assign _02629_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101101;
  assign _02630_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101100;
  assign _02631_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101011;
  assign _02632_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101010;
  assign _02633_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101001;
  assign _02634_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b101000;
  assign _02635_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100111;
  assign _02636_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100110;
  assign _02637_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100101;
  assign _02638_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100100;
  assign _02639_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100011;
  assign _02640_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100010;
  assign _02641_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100001;
  assign _02642_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 6'b100000;
  assign _02643_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11111;
  assign _02644_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11110;
  assign _02645_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11101;
  assign _02646_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11100;
  assign _02647_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11011;
  assign _02648_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11010;
  assign _02649_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11001;
  assign _02650_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b11000;
  assign _02651_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10111;
  assign _02652_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10110;
  assign _02653_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10101;
  assign _02654_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10100;
  assign _02655_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10011;
  assign _02656_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10010;
  assign _02657_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10001;
  assign _02658_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 5'b10000;
  assign _02659_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1111;
  assign _02660_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1110;
  assign _02661_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1101;
  assign _02662_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1100;
  assign _02663_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1011;
  assign _02664_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1010;
  assign _02665_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1001;
  assign _02666_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 4'b1000;
  assign _02667_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 3'b111;
  assign _02668_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 3'b110;
  assign _02669_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 3'b101;
  assign _02670_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 3'b100;
  assign _02671_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 2'b11;
  assign _02672_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 2'b10;
  assign _02673_ = vec_sum_112_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11115" *) 1'b1;
  function [7:0] _12080_;
    input [7:0] a;
    input [895:0] b;
    input [111:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *)
    (* parallel_case *)
    casez (s)
      112'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12080_ = b[7:0];
      112'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12080_ = b[15:8];
      112'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12080_ = b[23:16];
      112'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12080_ = b[31:24];
      112'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12080_ = b[39:32];
      112'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12080_ = b[47:40];
      112'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12080_ = b[55:48];
      112'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12080_ = b[63:56];
      112'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12080_ = b[71:64];
      112'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12080_ = b[79:72];
      112'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12080_ = b[87:80];
      112'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12080_ = b[95:88];
      112'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12080_ = b[103:96];
      112'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12080_ = b[111:104];
      112'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12080_ = b[119:112];
      112'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12080_ = b[127:120];
      112'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12080_ = b[135:128];
      112'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12080_ = b[143:136];
      112'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12080_ = b[151:144];
      112'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12080_ = b[159:152];
      112'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12080_ = b[167:160];
      112'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12080_ = b[175:168];
      112'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12080_ = b[183:176];
      112'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12080_ = b[191:184];
      112'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12080_ = b[199:192];
      112'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12080_ = b[207:200];
      112'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12080_ = b[215:208];
      112'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12080_ = b[223:216];
      112'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12080_ = b[231:224];
      112'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12080_ = b[239:232];
      112'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12080_ = b[247:240];
      112'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12080_ = b[255:248];
      112'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12080_ = b[263:256];
      112'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12080_ = b[271:264];
      112'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12080_ = b[279:272];
      112'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12080_ = b[287:280];
      112'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12080_ = b[295:288];
      112'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12080_ = b[303:296];
      112'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12080_ = b[311:304];
      112'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12080_ = b[319:312];
      112'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12080_ = b[327:320];
      112'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12080_ = b[335:328];
      112'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12080_ = b[343:336];
      112'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12080_ = b[351:344];
      112'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12080_ = b[359:352];
      112'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12080_ = b[367:360];
      112'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12080_ = b[375:368];
      112'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12080_ = b[383:376];
      112'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12080_ = b[391:384];
      112'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12080_ = b[399:392];
      112'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12080_ = b[407:400];
      112'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12080_ = b[415:408];
      112'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12080_ = b[423:416];
      112'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12080_ = b[431:424];
      112'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12080_ = b[439:432];
      112'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12080_ = b[447:440];
      112'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12080_ = b[455:448];
      112'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12080_ = b[463:456];
      112'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12080_ = b[471:464];
      112'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12080_ = b[479:472];
      112'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12080_ = b[487:480];
      112'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12080_ = b[495:488];
      112'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12080_ = b[503:496];
      112'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12080_ = b[511:504];
      112'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12080_ = b[519:512];
      112'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12080_ = b[527:520];
      112'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12080_ = b[535:528];
      112'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12080_ = b[543:536];
      112'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12080_ = b[551:544];
      112'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12080_ = b[559:552];
      112'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12080_ = b[567:560];
      112'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12080_ = b[575:568];
      112'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12080_ = b[583:576];
      112'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12080_ = b[591:584];
      112'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12080_ = b[599:592];
      112'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12080_ = b[607:600];
      112'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[615:608];
      112'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[623:616];
      112'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[631:624];
      112'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[639:632];
      112'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[647:640];
      112'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[655:648];
      112'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[663:656];
      112'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[671:664];
      112'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[679:672];
      112'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[687:680];
      112'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[695:688];
      112'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[703:696];
      112'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[711:704];
      112'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[719:712];
      112'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[727:720];
      112'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[735:728];
      112'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[743:736];
      112'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[751:744];
      112'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[759:752];
      112'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[767:760];
      112'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[775:768];
      112'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[783:776];
      112'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[791:784];
      112'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[799:792];
      112'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[807:800];
      112'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[815:808];
      112'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[823:816];
      112'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[831:824];
      112'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[839:832];
      112'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[847:840];
      112'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[855:848];
      112'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[863:856];
      112'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[871:864];
      112'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[879:872];
      112'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[887:880];
      112'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12080_ = b[895:888];
      default:
        _12080_ = a;
    endcase
  endfunction
  assign vec_data_111 = _12080_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880], data_d1[895:888] }, { _02785_, _02784_, _02783_, _02782_, _02781_, _02780_, _02779_, _02778_, _02777_, _02776_, _02775_, _02774_, _02773_, _02772_, _02771_, _02770_, _02769_, _02768_, _02767_, _02766_, _02765_, _02764_, _02763_, _02762_, _02761_, _02760_, _02759_, _02758_, _02757_, _02756_, _02755_, _02754_, _02753_, _02752_, _02751_, _02750_, _02749_, _02748_, _02747_, _02746_, _02745_, _02744_, _02743_, _02742_, _02741_, _02740_, _02739_, _02738_, _02737_, _02736_, _02735_, _02734_, _02733_, _02732_, _02731_, _02730_, _02729_, _02728_, _02727_, _02726_, _02725_, _02724_, _02723_, _02722_, _02721_, _02720_, _02719_, _02718_, _02717_, _02716_, _02715_, _02714_, _02713_, _02712_, _02711_, _02710_, _02709_, _02708_, _02707_, _02706_, _02705_, _02704_, _02703_, _02702_, _02701_, _02700_, _02699_, _02698_, _02697_, _02696_, _02695_, _02694_, _02693_, _02692_, _02691_, _02690_, _02689_, _02688_, _02687_, _02686_, _02685_, _02684_, _02683_, _02682_, _02681_, _02680_, _02679_, _02678_, _02677_, _02676_, _02675_, _02674_ });
  assign _02674_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1110000;
  assign _02675_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101111;
  assign _02676_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101110;
  assign _02677_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101101;
  assign _02678_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101100;
  assign _02679_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101011;
  assign _02680_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101010;
  assign _02681_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101001;
  assign _02682_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1101000;
  assign _02683_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100111;
  assign _02684_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100110;
  assign _02685_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100101;
  assign _02686_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100100;
  assign _02687_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100011;
  assign _02688_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100010;
  assign _02689_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100001;
  assign _02690_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1100000;
  assign _02691_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011111;
  assign _02692_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011110;
  assign _02693_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011101;
  assign _02694_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011100;
  assign _02695_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011011;
  assign _02696_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011010;
  assign _02697_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011001;
  assign _02698_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1011000;
  assign _02699_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010111;
  assign _02700_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010110;
  assign _02701_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010101;
  assign _02702_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010100;
  assign _02703_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010011;
  assign _02704_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010010;
  assign _02705_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010001;
  assign _02706_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1010000;
  assign _02707_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001111;
  assign _02708_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001110;
  assign _02709_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001101;
  assign _02710_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001100;
  assign _02711_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001011;
  assign _02712_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001010;
  assign _02713_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001001;
  assign _02714_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1001000;
  assign _02715_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000111;
  assign _02716_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000110;
  assign _02717_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000101;
  assign _02718_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000100;
  assign _02719_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000011;
  assign _02720_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000010;
  assign _02721_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000001;
  assign _02722_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 7'b1000000;
  assign _02723_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111111;
  assign _02724_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111110;
  assign _02725_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111101;
  assign _02726_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111100;
  assign _02727_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111011;
  assign _02728_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111010;
  assign _02729_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111001;
  assign _02730_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b111000;
  assign _02731_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110111;
  assign _02732_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110110;
  assign _02733_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110101;
  assign _02734_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110100;
  assign _02735_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110011;
  assign _02736_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110010;
  assign _02737_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110001;
  assign _02738_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b110000;
  assign _02739_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101111;
  assign _02740_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101110;
  assign _02741_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101101;
  assign _02742_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101100;
  assign _02743_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101011;
  assign _02744_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101010;
  assign _02745_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101001;
  assign _02746_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b101000;
  assign _02747_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100111;
  assign _02748_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100110;
  assign _02749_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100101;
  assign _02750_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100100;
  assign _02751_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100011;
  assign _02752_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100010;
  assign _02753_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100001;
  assign _02754_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 6'b100000;
  assign _02755_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11111;
  assign _02756_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11110;
  assign _02757_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11101;
  assign _02758_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11100;
  assign _02759_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11011;
  assign _02760_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11010;
  assign _02761_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11001;
  assign _02762_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b11000;
  assign _02763_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10111;
  assign _02764_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10110;
  assign _02765_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10101;
  assign _02766_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10100;
  assign _02767_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10011;
  assign _02768_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10010;
  assign _02769_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10001;
  assign _02770_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 5'b10000;
  assign _02771_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1111;
  assign _02772_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1110;
  assign _02773_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1101;
  assign _02774_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1100;
  assign _02775_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1011;
  assign _02776_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1010;
  assign _02777_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1001;
  assign _02778_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 4'b1000;
  assign _02779_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 3'b111;
  assign _02780_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 3'b110;
  assign _02781_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:11000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 3'b101;
  assign _02782_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 3'b100;
  assign _02783_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 2'b11;
  assign _02784_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 2'b10;
  assign _02785_ = vec_sum_111_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10995" *) 1'b1;
  function [7:0] _12193_;
    input [7:0] a;
    input [887:0] b;
    input [110:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *)
    (* parallel_case *)
    casez (s)
      111'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12193_ = b[7:0];
      111'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12193_ = b[15:8];
      111'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12193_ = b[23:16];
      111'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12193_ = b[31:24];
      111'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12193_ = b[39:32];
      111'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12193_ = b[47:40];
      111'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12193_ = b[55:48];
      111'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12193_ = b[63:56];
      111'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12193_ = b[71:64];
      111'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12193_ = b[79:72];
      111'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12193_ = b[87:80];
      111'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12193_ = b[95:88];
      111'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12193_ = b[103:96];
      111'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12193_ = b[111:104];
      111'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12193_ = b[119:112];
      111'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12193_ = b[127:120];
      111'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12193_ = b[135:128];
      111'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12193_ = b[143:136];
      111'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12193_ = b[151:144];
      111'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12193_ = b[159:152];
      111'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12193_ = b[167:160];
      111'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12193_ = b[175:168];
      111'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12193_ = b[183:176];
      111'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12193_ = b[191:184];
      111'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12193_ = b[199:192];
      111'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12193_ = b[207:200];
      111'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12193_ = b[215:208];
      111'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12193_ = b[223:216];
      111'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12193_ = b[231:224];
      111'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12193_ = b[239:232];
      111'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12193_ = b[247:240];
      111'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12193_ = b[255:248];
      111'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12193_ = b[263:256];
      111'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12193_ = b[271:264];
      111'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12193_ = b[279:272];
      111'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12193_ = b[287:280];
      111'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12193_ = b[295:288];
      111'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12193_ = b[303:296];
      111'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12193_ = b[311:304];
      111'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12193_ = b[319:312];
      111'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12193_ = b[327:320];
      111'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12193_ = b[335:328];
      111'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12193_ = b[343:336];
      111'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12193_ = b[351:344];
      111'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12193_ = b[359:352];
      111'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12193_ = b[367:360];
      111'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12193_ = b[375:368];
      111'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12193_ = b[383:376];
      111'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12193_ = b[391:384];
      111'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12193_ = b[399:392];
      111'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12193_ = b[407:400];
      111'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12193_ = b[415:408];
      111'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12193_ = b[423:416];
      111'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12193_ = b[431:424];
      111'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12193_ = b[439:432];
      111'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12193_ = b[447:440];
      111'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12193_ = b[455:448];
      111'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12193_ = b[463:456];
      111'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12193_ = b[471:464];
      111'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12193_ = b[479:472];
      111'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12193_ = b[487:480];
      111'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12193_ = b[495:488];
      111'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12193_ = b[503:496];
      111'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12193_ = b[511:504];
      111'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12193_ = b[519:512];
      111'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12193_ = b[527:520];
      111'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12193_ = b[535:528];
      111'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12193_ = b[543:536];
      111'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12193_ = b[551:544];
      111'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12193_ = b[559:552];
      111'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12193_ = b[567:560];
      111'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12193_ = b[575:568];
      111'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12193_ = b[583:576];
      111'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12193_ = b[591:584];
      111'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12193_ = b[599:592];
      111'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12193_ = b[607:600];
      111'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[615:608];
      111'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[623:616];
      111'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[631:624];
      111'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[639:632];
      111'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[647:640];
      111'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[655:648];
      111'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[663:656];
      111'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[671:664];
      111'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[679:672];
      111'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[687:680];
      111'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[695:688];
      111'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[703:696];
      111'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[711:704];
      111'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[719:712];
      111'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[727:720];
      111'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[735:728];
      111'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[743:736];
      111'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[751:744];
      111'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[759:752];
      111'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[767:760];
      111'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[775:768];
      111'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[783:776];
      111'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[791:784];
      111'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[799:792];
      111'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[807:800];
      111'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[815:808];
      111'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[823:816];
      111'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[831:824];
      111'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[839:832];
      111'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[847:840];
      111'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[855:848];
      111'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[863:856];
      111'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[871:864];
      111'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[879:872];
      111'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12193_ = b[887:880];
      default:
        _12193_ = a;
    endcase
  endfunction
  assign vec_data_110 = _12193_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872], data_d1[887:880] }, { _02896_, _02895_, _02894_, _02893_, _02892_, _02891_, _02890_, _02889_, _02888_, _02887_, _02886_, _02885_, _02884_, _02883_, _02882_, _02881_, _02880_, _02879_, _02878_, _02877_, _02876_, _02875_, _02874_, _02873_, _02872_, _02871_, _02870_, _02869_, _02868_, _02867_, _02866_, _02865_, _02864_, _02863_, _02862_, _02861_, _02860_, _02859_, _02858_, _02857_, _02856_, _02855_, _02854_, _02853_, _02852_, _02851_, _02850_, _02849_, _02848_, _02847_, _02846_, _02845_, _02844_, _02843_, _02842_, _02841_, _02840_, _02839_, _02838_, _02837_, _02836_, _02835_, _02834_, _02833_, _02832_, _02831_, _02830_, _02829_, _02828_, _02827_, _02826_, _02825_, _02824_, _02823_, _02822_, _02821_, _02820_, _02819_, _02818_, _02817_, _02816_, _02815_, _02814_, _02813_, _02812_, _02811_, _02810_, _02809_, _02808_, _02807_, _02806_, _02805_, _02804_, _02803_, _02802_, _02801_, _02800_, _02799_, _02798_, _02797_, _02796_, _02795_, _02794_, _02793_, _02792_, _02791_, _02790_, _02789_, _02788_, _02787_, _02786_ });
  assign _02786_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101111;
  assign _02787_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101110;
  assign _02788_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101101;
  assign _02789_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101100;
  assign _02790_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101011;
  assign _02791_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101010;
  assign _02792_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101001;
  assign _02793_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1101000;
  assign _02794_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100111;
  assign _02795_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100110;
  assign _02796_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100101;
  assign _02797_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100100;
  assign _02798_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100011;
  assign _02799_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100010;
  assign _02800_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100001;
  assign _02801_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1100000;
  assign _02802_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011111;
  assign _02803_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011110;
  assign _02804_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011101;
  assign _02805_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011100;
  assign _02806_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011011;
  assign _02807_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011010;
  assign _02808_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011001;
  assign _02809_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1011000;
  assign _02810_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010111;
  assign _02811_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010110;
  assign _02812_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010101;
  assign _02813_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010100;
  assign _02814_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010011;
  assign _02815_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010010;
  assign _02816_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010001;
  assign _02817_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1010000;
  assign _02818_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001111;
  assign _02819_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001110;
  assign _02820_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001101;
  assign _02821_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001100;
  assign _02822_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001011;
  assign _02823_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001010;
  assign _02824_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001001;
  assign _02825_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1001000;
  assign _02826_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000111;
  assign _02827_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000110;
  assign _02828_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000101;
  assign _02829_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000100;
  assign _02830_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000011;
  assign _02831_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000010;
  assign _02832_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000001;
  assign _02833_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 7'b1000000;
  assign _02834_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111111;
  assign _02835_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111110;
  assign _02836_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111101;
  assign _02837_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111100;
  assign _02838_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111011;
  assign _02839_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111010;
  assign _02840_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111001;
  assign _02841_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b111000;
  assign _02842_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110111;
  assign _02843_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110110;
  assign _02844_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110101;
  assign _02845_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110100;
  assign _02846_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110011;
  assign _02847_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110010;
  assign _02848_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110001;
  assign _02849_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b110000;
  assign _02850_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101111;
  assign _02851_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101110;
  assign _02852_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101101;
  assign _02853_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101100;
  assign _02854_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101011;
  assign _02855_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101010;
  assign _02856_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101001;
  assign _02857_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b101000;
  assign _02858_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100111;
  assign _02859_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100110;
  assign _02860_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100101;
  assign _02861_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100100;
  assign _02862_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100011;
  assign _02863_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100010;
  assign _02864_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100001;
  assign _02865_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 6'b100000;
  assign _02866_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11111;
  assign _02867_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11110;
  assign _02868_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11101;
  assign _02869_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11100;
  assign _02870_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11011;
  assign _02871_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11010;
  assign _02872_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11001;
  assign _02873_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b11000;
  assign _02874_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10111;
  assign _02875_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10110;
  assign _02876_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10101;
  assign _02877_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10100;
  assign _02878_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10011;
  assign _02879_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10010;
  assign _02880_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10001;
  assign _02881_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 5'b10000;
  assign _02882_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1111;
  assign _02883_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1110;
  assign _02884_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1101;
  assign _02885_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1100;
  assign _02886_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1011;
  assign _02887_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1010;
  assign _02888_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1001;
  assign _02889_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 4'b1000;
  assign _02890_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 3'b111;
  assign _02891_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 3'b110;
  assign _02892_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 3'b101;
  assign _02893_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 3'b100;
  assign _02894_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 2'b11;
  assign _02895_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 2'b10;
  assign _02896_ = vec_sum_110_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10876" *) 1'b1;
  function [7:0] _12305_;
    input [7:0] a;
    input [879:0] b;
    input [109:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *)
    (* parallel_case *)
    casez (s)
      110'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12305_ = b[7:0];
      110'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12305_ = b[15:8];
      110'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12305_ = b[23:16];
      110'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12305_ = b[31:24];
      110'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12305_ = b[39:32];
      110'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12305_ = b[47:40];
      110'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12305_ = b[55:48];
      110'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12305_ = b[63:56];
      110'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12305_ = b[71:64];
      110'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12305_ = b[79:72];
      110'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12305_ = b[87:80];
      110'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12305_ = b[95:88];
      110'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12305_ = b[103:96];
      110'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12305_ = b[111:104];
      110'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12305_ = b[119:112];
      110'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12305_ = b[127:120];
      110'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12305_ = b[135:128];
      110'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12305_ = b[143:136];
      110'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12305_ = b[151:144];
      110'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12305_ = b[159:152];
      110'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12305_ = b[167:160];
      110'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12305_ = b[175:168];
      110'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12305_ = b[183:176];
      110'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12305_ = b[191:184];
      110'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12305_ = b[199:192];
      110'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12305_ = b[207:200];
      110'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12305_ = b[215:208];
      110'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12305_ = b[223:216];
      110'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12305_ = b[231:224];
      110'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12305_ = b[239:232];
      110'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12305_ = b[247:240];
      110'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12305_ = b[255:248];
      110'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12305_ = b[263:256];
      110'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12305_ = b[271:264];
      110'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12305_ = b[279:272];
      110'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12305_ = b[287:280];
      110'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12305_ = b[295:288];
      110'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12305_ = b[303:296];
      110'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12305_ = b[311:304];
      110'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12305_ = b[319:312];
      110'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12305_ = b[327:320];
      110'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12305_ = b[335:328];
      110'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12305_ = b[343:336];
      110'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12305_ = b[351:344];
      110'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12305_ = b[359:352];
      110'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12305_ = b[367:360];
      110'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12305_ = b[375:368];
      110'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12305_ = b[383:376];
      110'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12305_ = b[391:384];
      110'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12305_ = b[399:392];
      110'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12305_ = b[407:400];
      110'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12305_ = b[415:408];
      110'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12305_ = b[423:416];
      110'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12305_ = b[431:424];
      110'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12305_ = b[439:432];
      110'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12305_ = b[447:440];
      110'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12305_ = b[455:448];
      110'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12305_ = b[463:456];
      110'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12305_ = b[471:464];
      110'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12305_ = b[479:472];
      110'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12305_ = b[487:480];
      110'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12305_ = b[495:488];
      110'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12305_ = b[503:496];
      110'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12305_ = b[511:504];
      110'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12305_ = b[519:512];
      110'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12305_ = b[527:520];
      110'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12305_ = b[535:528];
      110'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12305_ = b[543:536];
      110'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12305_ = b[551:544];
      110'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12305_ = b[559:552];
      110'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12305_ = b[567:560];
      110'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12305_ = b[575:568];
      110'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12305_ = b[583:576];
      110'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12305_ = b[591:584];
      110'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12305_ = b[599:592];
      110'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12305_ = b[607:600];
      110'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[615:608];
      110'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[623:616];
      110'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[631:624];
      110'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[639:632];
      110'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[647:640];
      110'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[655:648];
      110'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[663:656];
      110'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[671:664];
      110'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[679:672];
      110'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[687:680];
      110'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[695:688];
      110'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[703:696];
      110'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[711:704];
      110'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[719:712];
      110'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[727:720];
      110'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[735:728];
      110'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[743:736];
      110'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[751:744];
      110'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[759:752];
      110'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[767:760];
      110'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[775:768];
      110'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[783:776];
      110'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[791:784];
      110'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[799:792];
      110'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[807:800];
      110'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[815:808];
      110'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[823:816];
      110'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[831:824];
      110'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[839:832];
      110'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[847:840];
      110'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[855:848];
      110'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[863:856];
      110'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[871:864];
      110'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12305_ = b[879:872];
      default:
        _12305_ = a;
    endcase
  endfunction
  assign vec_data_109 = _12305_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864], data_d1[879:872] }, { _03006_, _03005_, _03004_, _03003_, _03002_, _03001_, _03000_, _02999_, _02998_, _02997_, _02996_, _02995_, _02994_, _02993_, _02992_, _02991_, _02990_, _02989_, _02988_, _02987_, _02986_, _02985_, _02984_, _02983_, _02982_, _02981_, _02980_, _02979_, _02978_, _02977_, _02976_, _02975_, _02974_, _02973_, _02972_, _02971_, _02970_, _02969_, _02968_, _02967_, _02966_, _02965_, _02964_, _02963_, _02962_, _02961_, _02960_, _02959_, _02958_, _02957_, _02956_, _02955_, _02954_, _02953_, _02952_, _02951_, _02950_, _02949_, _02948_, _02947_, _02946_, _02945_, _02944_, _02943_, _02942_, _02941_, _02940_, _02939_, _02938_, _02937_, _02936_, _02935_, _02934_, _02933_, _02932_, _02931_, _02930_, _02929_, _02928_, _02927_, _02926_, _02925_, _02924_, _02923_, _02922_, _02921_, _02920_, _02919_, _02918_, _02917_, _02916_, _02915_, _02914_, _02913_, _02912_, _02911_, _02910_, _02909_, _02908_, _02907_, _02906_, _02905_, _02904_, _02903_, _02902_, _02901_, _02900_, _02899_, _02898_, _02897_ });
  assign _02897_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101110;
  assign _02898_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101101;
  assign _02899_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101100;
  assign _02900_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101011;
  assign _02901_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101010;
  assign _02902_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101001;
  assign _02903_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1101000;
  assign _02904_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100111;
  assign _02905_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100110;
  assign _02906_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100101;
  assign _02907_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100100;
  assign _02908_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100011;
  assign _02909_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100010;
  assign _02910_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100001;
  assign _02911_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1100000;
  assign _02912_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011111;
  assign _02913_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011110;
  assign _02914_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011101;
  assign _02915_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011100;
  assign _02916_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011011;
  assign _02917_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011010;
  assign _02918_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011001;
  assign _02919_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1011000;
  assign _02920_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010111;
  assign _02921_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010110;
  assign _02922_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010101;
  assign _02923_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010100;
  assign _02924_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010011;
  assign _02925_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010010;
  assign _02926_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010001;
  assign _02927_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1010000;
  assign _02928_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001111;
  assign _02929_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001110;
  assign _02930_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001101;
  assign _02931_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001100;
  assign _02932_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001011;
  assign _02933_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001010;
  assign _02934_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001001;
  assign _02935_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1001000;
  assign _02936_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000111;
  assign _02937_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000110;
  assign _02938_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000101;
  assign _02939_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000100;
  assign _02940_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000011;
  assign _02941_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000010;
  assign _02942_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000001;
  assign _02943_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 7'b1000000;
  assign _02944_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111111;
  assign _02945_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111110;
  assign _02946_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111101;
  assign _02947_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111100;
  assign _02948_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111011;
  assign _02949_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111010;
  assign _02950_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111001;
  assign _02951_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b111000;
  assign _02952_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110111;
  assign _02953_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110110;
  assign _02954_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110101;
  assign _02955_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110100;
  assign _02956_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110011;
  assign _02957_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110010;
  assign _02958_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110001;
  assign _02959_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b110000;
  assign _02960_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101111;
  assign _02961_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101110;
  assign _02962_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101101;
  assign _02963_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101100;
  assign _02964_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101011;
  assign _02965_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101010;
  assign _02966_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101001;
  assign _02967_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b101000;
  assign _02968_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100111;
  assign _02969_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100110;
  assign _02970_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100101;
  assign _02971_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100100;
  assign _02972_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100011;
  assign _02973_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100010;
  assign _02974_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100001;
  assign _02975_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 6'b100000;
  assign _02976_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11111;
  assign _02977_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11110;
  assign _02978_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11101;
  assign _02979_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11100;
  assign _02980_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11011;
  assign _02981_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11010;
  assign _02982_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11001;
  assign _02983_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b11000;
  assign _02984_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10111;
  assign _02985_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10110;
  assign _02986_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10101;
  assign _02987_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10100;
  assign _02988_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10011;
  assign _02989_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10010;
  assign _02990_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10001;
  assign _02991_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 5'b10000;
  assign _02992_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1111;
  assign _02993_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1110;
  assign _02994_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1101;
  assign _02995_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1100;
  assign _02996_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1011;
  assign _02997_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1010;
  assign _02998_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1001;
  assign _02999_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 4'b1000;
  assign _03000_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 3'b111;
  assign _03001_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 3'b110;
  assign _03002_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 3'b101;
  assign _03003_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 3'b100;
  assign _03004_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 2'b11;
  assign _03005_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 2'b10;
  assign _03006_ = vec_sum_109_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10758" *) 1'b1;
  function [7:0] _12416_;
    input [7:0] a;
    input [871:0] b;
    input [108:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *)
    (* parallel_case *)
    casez (s)
      109'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12416_ = b[7:0];
      109'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12416_ = b[15:8];
      109'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12416_ = b[23:16];
      109'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12416_ = b[31:24];
      109'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12416_ = b[39:32];
      109'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12416_ = b[47:40];
      109'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12416_ = b[55:48];
      109'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12416_ = b[63:56];
      109'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12416_ = b[71:64];
      109'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12416_ = b[79:72];
      109'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12416_ = b[87:80];
      109'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12416_ = b[95:88];
      109'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12416_ = b[103:96];
      109'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12416_ = b[111:104];
      109'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12416_ = b[119:112];
      109'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12416_ = b[127:120];
      109'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12416_ = b[135:128];
      109'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12416_ = b[143:136];
      109'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12416_ = b[151:144];
      109'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12416_ = b[159:152];
      109'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12416_ = b[167:160];
      109'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12416_ = b[175:168];
      109'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12416_ = b[183:176];
      109'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12416_ = b[191:184];
      109'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12416_ = b[199:192];
      109'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12416_ = b[207:200];
      109'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12416_ = b[215:208];
      109'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12416_ = b[223:216];
      109'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12416_ = b[231:224];
      109'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12416_ = b[239:232];
      109'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12416_ = b[247:240];
      109'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12416_ = b[255:248];
      109'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12416_ = b[263:256];
      109'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12416_ = b[271:264];
      109'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12416_ = b[279:272];
      109'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12416_ = b[287:280];
      109'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12416_ = b[295:288];
      109'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12416_ = b[303:296];
      109'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12416_ = b[311:304];
      109'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12416_ = b[319:312];
      109'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12416_ = b[327:320];
      109'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12416_ = b[335:328];
      109'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12416_ = b[343:336];
      109'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12416_ = b[351:344];
      109'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12416_ = b[359:352];
      109'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12416_ = b[367:360];
      109'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12416_ = b[375:368];
      109'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12416_ = b[383:376];
      109'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12416_ = b[391:384];
      109'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12416_ = b[399:392];
      109'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12416_ = b[407:400];
      109'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12416_ = b[415:408];
      109'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12416_ = b[423:416];
      109'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12416_ = b[431:424];
      109'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12416_ = b[439:432];
      109'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12416_ = b[447:440];
      109'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12416_ = b[455:448];
      109'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12416_ = b[463:456];
      109'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12416_ = b[471:464];
      109'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12416_ = b[479:472];
      109'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12416_ = b[487:480];
      109'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12416_ = b[495:488];
      109'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12416_ = b[503:496];
      109'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12416_ = b[511:504];
      109'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12416_ = b[519:512];
      109'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12416_ = b[527:520];
      109'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12416_ = b[535:528];
      109'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12416_ = b[543:536];
      109'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12416_ = b[551:544];
      109'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12416_ = b[559:552];
      109'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12416_ = b[567:560];
      109'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12416_ = b[575:568];
      109'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12416_ = b[583:576];
      109'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12416_ = b[591:584];
      109'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12416_ = b[599:592];
      109'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12416_ = b[607:600];
      109'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[615:608];
      109'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[623:616];
      109'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[631:624];
      109'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[639:632];
      109'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[647:640];
      109'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[655:648];
      109'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[663:656];
      109'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[671:664];
      109'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[679:672];
      109'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[687:680];
      109'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[695:688];
      109'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[703:696];
      109'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[711:704];
      109'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[719:712];
      109'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[727:720];
      109'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[735:728];
      109'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[743:736];
      109'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[751:744];
      109'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[759:752];
      109'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[767:760];
      109'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[775:768];
      109'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[783:776];
      109'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[791:784];
      109'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[799:792];
      109'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[807:800];
      109'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[815:808];
      109'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[823:816];
      109'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[831:824];
      109'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[839:832];
      109'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[847:840];
      109'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[855:848];
      109'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[863:856];
      109'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12416_ = b[871:864];
      default:
        _12416_ = a;
    endcase
  endfunction
  assign vec_data_108 = _12416_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856], data_d1[871:864] }, { _03115_, _03114_, _03113_, _03112_, _03111_, _03110_, _03109_, _03108_, _03107_, _03106_, _03105_, _03104_, _03103_, _03102_, _03101_, _03100_, _03099_, _03098_, _03097_, _03096_, _03095_, _03094_, _03093_, _03092_, _03091_, _03090_, _03089_, _03088_, _03087_, _03086_, _03085_, _03084_, _03083_, _03082_, _03081_, _03080_, _03079_, _03078_, _03077_, _03076_, _03075_, _03074_, _03073_, _03072_, _03071_, _03070_, _03069_, _03068_, _03067_, _03066_, _03065_, _03064_, _03063_, _03062_, _03061_, _03060_, _03059_, _03058_, _03057_, _03056_, _03055_, _03054_, _03053_, _03052_, _03051_, _03050_, _03049_, _03048_, _03047_, _03046_, _03045_, _03044_, _03043_, _03042_, _03041_, _03040_, _03039_, _03038_, _03037_, _03036_, _03035_, _03034_, _03033_, _03032_, _03031_, _03030_, _03029_, _03028_, _03027_, _03026_, _03025_, _03024_, _03023_, _03022_, _03021_, _03020_, _03019_, _03018_, _03017_, _03016_, _03015_, _03014_, _03013_, _03012_, _03011_, _03010_, _03009_, _03008_, _03007_ });
  assign _03007_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101101;
  assign _03008_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101100;
  assign _03009_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101011;
  assign _03010_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101010;
  assign _03011_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101001;
  assign _03012_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1101000;
  assign _03013_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100111;
  assign _03014_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100110;
  assign _03015_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100101;
  assign _03016_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100100;
  assign _03017_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100011;
  assign _03018_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100010;
  assign _03019_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100001;
  assign _03020_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1100000;
  assign _03021_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011111;
  assign _03022_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011110;
  assign _03023_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011101;
  assign _03024_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011100;
  assign _03025_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011011;
  assign _03026_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011010;
  assign _03027_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011001;
  assign _03028_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1011000;
  assign _03029_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010111;
  assign _03030_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010110;
  assign _03031_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010101;
  assign _03032_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010100;
  assign _03033_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010011;
  assign _03034_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010010;
  assign _03035_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010001;
  assign _03036_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1010000;
  assign _03037_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001111;
  assign _03038_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001110;
  assign _03039_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001101;
  assign _03040_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001100;
  assign _03041_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001011;
  assign _03042_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001010;
  assign _03043_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001001;
  assign _03044_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1001000;
  assign _03045_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000111;
  assign _03046_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000110;
  assign _03047_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000101;
  assign _03048_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000100;
  assign _03049_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000011;
  assign _03050_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000010;
  assign _03051_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000001;
  assign _03052_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 7'b1000000;
  assign _03053_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111111;
  assign _03054_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111110;
  assign _03055_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111101;
  assign _03056_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111100;
  assign _03057_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111011;
  assign _03058_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111010;
  assign _03059_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111001;
  assign _03060_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b111000;
  assign _03061_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110111;
  assign _03062_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110110;
  assign _03063_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110101;
  assign _03064_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110100;
  assign _03065_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110011;
  assign _03066_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110010;
  assign _03067_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110001;
  assign _03068_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b110000;
  assign _03069_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101111;
  assign _03070_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101110;
  assign _03071_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101101;
  assign _03072_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101100;
  assign _03073_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101011;
  assign _03074_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101010;
  assign _03075_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101001;
  assign _03076_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b101000;
  assign _03077_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100111;
  assign _03078_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100110;
  assign _03079_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100101;
  assign _03080_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100100;
  assign _03081_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100011;
  assign _03082_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100010;
  assign _03083_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100001;
  assign _03084_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 6'b100000;
  assign _03085_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11111;
  assign _03086_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11110;
  assign _03087_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11101;
  assign _03088_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11100;
  assign _03089_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11011;
  assign _03090_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11010;
  assign _03091_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11001;
  assign _03092_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b11000;
  assign _03093_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10111;
  assign _03094_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10110;
  assign _03095_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10101;
  assign _03096_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10100;
  assign _03097_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10011;
  assign _03098_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10010;
  assign _03099_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10001;
  assign _03100_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 5'b10000;
  assign _03101_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1111;
  assign _03102_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1110;
  assign _03103_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1101;
  assign _03104_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1100;
  assign _03105_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1011;
  assign _03106_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1010;
  assign _03107_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1001;
  assign _03108_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 4'b1000;
  assign _03109_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 3'b111;
  assign _03110_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 3'b110;
  assign _03111_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 3'b101;
  assign _03112_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 3'b100;
  assign _03113_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 2'b11;
  assign _03114_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 2'b10;
  assign _03115_ = vec_sum_108_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10641" *) 1'b1;
  function [7:0] _12526_;
    input [7:0] a;
    input [863:0] b;
    input [107:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *)
    (* parallel_case *)
    casez (s)
      108'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12526_ = b[7:0];
      108'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12526_ = b[15:8];
      108'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12526_ = b[23:16];
      108'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12526_ = b[31:24];
      108'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12526_ = b[39:32];
      108'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12526_ = b[47:40];
      108'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12526_ = b[55:48];
      108'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12526_ = b[63:56];
      108'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12526_ = b[71:64];
      108'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12526_ = b[79:72];
      108'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12526_ = b[87:80];
      108'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12526_ = b[95:88];
      108'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12526_ = b[103:96];
      108'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12526_ = b[111:104];
      108'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12526_ = b[119:112];
      108'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12526_ = b[127:120];
      108'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12526_ = b[135:128];
      108'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12526_ = b[143:136];
      108'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12526_ = b[151:144];
      108'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12526_ = b[159:152];
      108'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12526_ = b[167:160];
      108'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12526_ = b[175:168];
      108'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12526_ = b[183:176];
      108'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12526_ = b[191:184];
      108'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12526_ = b[199:192];
      108'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12526_ = b[207:200];
      108'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12526_ = b[215:208];
      108'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12526_ = b[223:216];
      108'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12526_ = b[231:224];
      108'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12526_ = b[239:232];
      108'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12526_ = b[247:240];
      108'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12526_ = b[255:248];
      108'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12526_ = b[263:256];
      108'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12526_ = b[271:264];
      108'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12526_ = b[279:272];
      108'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12526_ = b[287:280];
      108'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12526_ = b[295:288];
      108'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12526_ = b[303:296];
      108'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12526_ = b[311:304];
      108'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12526_ = b[319:312];
      108'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12526_ = b[327:320];
      108'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12526_ = b[335:328];
      108'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12526_ = b[343:336];
      108'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12526_ = b[351:344];
      108'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12526_ = b[359:352];
      108'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12526_ = b[367:360];
      108'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12526_ = b[375:368];
      108'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12526_ = b[383:376];
      108'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12526_ = b[391:384];
      108'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12526_ = b[399:392];
      108'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12526_ = b[407:400];
      108'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12526_ = b[415:408];
      108'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12526_ = b[423:416];
      108'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12526_ = b[431:424];
      108'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12526_ = b[439:432];
      108'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12526_ = b[447:440];
      108'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12526_ = b[455:448];
      108'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12526_ = b[463:456];
      108'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12526_ = b[471:464];
      108'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12526_ = b[479:472];
      108'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12526_ = b[487:480];
      108'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12526_ = b[495:488];
      108'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12526_ = b[503:496];
      108'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12526_ = b[511:504];
      108'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12526_ = b[519:512];
      108'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12526_ = b[527:520];
      108'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12526_ = b[535:528];
      108'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12526_ = b[543:536];
      108'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12526_ = b[551:544];
      108'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12526_ = b[559:552];
      108'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12526_ = b[567:560];
      108'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12526_ = b[575:568];
      108'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12526_ = b[583:576];
      108'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12526_ = b[591:584];
      108'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12526_ = b[599:592];
      108'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12526_ = b[607:600];
      108'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[615:608];
      108'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[623:616];
      108'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[631:624];
      108'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[639:632];
      108'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[647:640];
      108'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[655:648];
      108'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[663:656];
      108'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[671:664];
      108'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[679:672];
      108'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[687:680];
      108'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[695:688];
      108'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[703:696];
      108'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[711:704];
      108'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[719:712];
      108'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[727:720];
      108'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[735:728];
      108'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[743:736];
      108'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[751:744];
      108'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[759:752];
      108'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[767:760];
      108'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[775:768];
      108'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[783:776];
      108'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[791:784];
      108'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[799:792];
      108'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[807:800];
      108'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[815:808];
      108'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[823:816];
      108'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[831:824];
      108'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[839:832];
      108'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[847:840];
      108'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[855:848];
      108'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12526_ = b[863:856];
      default:
        _12526_ = a;
    endcase
  endfunction
  assign vec_data_107 = _12526_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848], data_d1[863:856] }, { _03223_, _03222_, _03221_, _03220_, _03219_, _03218_, _03217_, _03216_, _03215_, _03214_, _03213_, _03212_, _03211_, _03210_, _03209_, _03208_, _03207_, _03206_, _03205_, _03204_, _03203_, _03202_, _03201_, _03200_, _03199_, _03198_, _03197_, _03196_, _03195_, _03194_, _03193_, _03192_, _03191_, _03190_, _03189_, _03188_, _03187_, _03186_, _03185_, _03184_, _03183_, _03182_, _03181_, _03180_, _03179_, _03178_, _03177_, _03176_, _03175_, _03174_, _03173_, _03172_, _03171_, _03170_, _03169_, _03168_, _03167_, _03166_, _03165_, _03164_, _03163_, _03162_, _03161_, _03160_, _03159_, _03158_, _03157_, _03156_, _03155_, _03154_, _03153_, _03152_, _03151_, _03150_, _03149_, _03148_, _03147_, _03146_, _03145_, _03144_, _03143_, _03142_, _03141_, _03140_, _03139_, _03138_, _03137_, _03136_, _03135_, _03134_, _03133_, _03132_, _03131_, _03130_, _03129_, _03128_, _03127_, _03126_, _03125_, _03124_, _03123_, _03122_, _03121_, _03120_, _03119_, _03118_, _03117_, _03116_ });
  assign _03116_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1101100;
  assign _03117_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1101011;
  assign _03118_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1101010;
  assign _03119_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10630|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1101001;
  assign _03120_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10629|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1101000;
  assign _03121_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10628|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100111;
  assign _03122_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100110;
  assign _03123_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100101;
  assign _03124_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100100;
  assign _03125_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100011;
  assign _03126_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100010;
  assign _03127_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100001;
  assign _03128_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1100000;
  assign _03129_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011111;
  assign _03130_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011110;
  assign _03131_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011101;
  assign _03132_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011100;
  assign _03133_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011011;
  assign _03134_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011010;
  assign _03135_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011001;
  assign _03136_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1011000;
  assign _03137_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010111;
  assign _03138_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010110;
  assign _03139_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010101;
  assign _03140_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010100;
  assign _03141_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010011;
  assign _03142_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010010;
  assign _03143_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010001;
  assign _03144_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1010000;
  assign _03145_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001111;
  assign _03146_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001110;
  assign _03147_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001101;
  assign _03148_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001100;
  assign _03149_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001011;
  assign _03150_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001010;
  assign _03151_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001001;
  assign _03152_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1001000;
  assign _03153_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000111;
  assign _03154_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000110;
  assign _03155_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000101;
  assign _03156_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000100;
  assign _03157_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000011;
  assign _03158_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000010;
  assign _03159_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000001;
  assign _03160_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 7'b1000000;
  assign _03161_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111111;
  assign _03162_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111110;
  assign _03163_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111101;
  assign _03164_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111100;
  assign _03165_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111011;
  assign _03166_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111010;
  assign _03167_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111001;
  assign _03168_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b111000;
  assign _03169_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110111;
  assign _03170_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110110;
  assign _03171_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110101;
  assign _03172_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110100;
  assign _03173_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110011;
  assign _03174_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110010;
  assign _03175_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110001;
  assign _03176_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b110000;
  assign _03177_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101111;
  assign _03178_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101110;
  assign _03179_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101101;
  assign _03180_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101100;
  assign _03181_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101011;
  assign _03182_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101010;
  assign _03183_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101001;
  assign _03184_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b101000;
  assign _03185_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100111;
  assign _03186_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100110;
  assign _03187_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100101;
  assign _03188_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100100;
  assign _03189_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100011;
  assign _03190_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100010;
  assign _03191_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100001;
  assign _03192_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 6'b100000;
  assign _03193_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11111;
  assign _03194_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11110;
  assign _03195_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11101;
  assign _03196_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11100;
  assign _03197_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11011;
  assign _03198_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11010;
  assign _03199_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11001;
  assign _03200_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b11000;
  assign _03201_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10111;
  assign _03202_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10110;
  assign _03203_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10101;
  assign _03204_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10100;
  assign _03205_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10011;
  assign _03206_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10010;
  assign _03207_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10001;
  assign _03208_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 5'b10000;
  assign _03209_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1111;
  assign _03210_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1110;
  assign _03211_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1101;
  assign _03212_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1100;
  assign _03213_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1011;
  assign _03214_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1010;
  assign _03215_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1001;
  assign _03216_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 4'b1000;
  assign _03217_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 3'b111;
  assign _03218_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 3'b110;
  assign _03219_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 3'b101;
  assign _03220_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 3'b100;
  assign _03221_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 2'b11;
  assign _03222_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 2'b10;
  assign _03223_ = vec_sum_107_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10525" *) 1'b1;
  function [7:0] _12635_;
    input [7:0] a;
    input [855:0] b;
    input [106:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *)
    (* parallel_case *)
    casez (s)
      107'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12635_ = b[7:0];
      107'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12635_ = b[15:8];
      107'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12635_ = b[23:16];
      107'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12635_ = b[31:24];
      107'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12635_ = b[39:32];
      107'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12635_ = b[47:40];
      107'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12635_ = b[55:48];
      107'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12635_ = b[63:56];
      107'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12635_ = b[71:64];
      107'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12635_ = b[79:72];
      107'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12635_ = b[87:80];
      107'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12635_ = b[95:88];
      107'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12635_ = b[103:96];
      107'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12635_ = b[111:104];
      107'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12635_ = b[119:112];
      107'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12635_ = b[127:120];
      107'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12635_ = b[135:128];
      107'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12635_ = b[143:136];
      107'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12635_ = b[151:144];
      107'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12635_ = b[159:152];
      107'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12635_ = b[167:160];
      107'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12635_ = b[175:168];
      107'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12635_ = b[183:176];
      107'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12635_ = b[191:184];
      107'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12635_ = b[199:192];
      107'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12635_ = b[207:200];
      107'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12635_ = b[215:208];
      107'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12635_ = b[223:216];
      107'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12635_ = b[231:224];
      107'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12635_ = b[239:232];
      107'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12635_ = b[247:240];
      107'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12635_ = b[255:248];
      107'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12635_ = b[263:256];
      107'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12635_ = b[271:264];
      107'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12635_ = b[279:272];
      107'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12635_ = b[287:280];
      107'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12635_ = b[295:288];
      107'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12635_ = b[303:296];
      107'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12635_ = b[311:304];
      107'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12635_ = b[319:312];
      107'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12635_ = b[327:320];
      107'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12635_ = b[335:328];
      107'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12635_ = b[343:336];
      107'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12635_ = b[351:344];
      107'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12635_ = b[359:352];
      107'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12635_ = b[367:360];
      107'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12635_ = b[375:368];
      107'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12635_ = b[383:376];
      107'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12635_ = b[391:384];
      107'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12635_ = b[399:392];
      107'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12635_ = b[407:400];
      107'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12635_ = b[415:408];
      107'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12635_ = b[423:416];
      107'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12635_ = b[431:424];
      107'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12635_ = b[439:432];
      107'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12635_ = b[447:440];
      107'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12635_ = b[455:448];
      107'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12635_ = b[463:456];
      107'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12635_ = b[471:464];
      107'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12635_ = b[479:472];
      107'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12635_ = b[487:480];
      107'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12635_ = b[495:488];
      107'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12635_ = b[503:496];
      107'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12635_ = b[511:504];
      107'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12635_ = b[519:512];
      107'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12635_ = b[527:520];
      107'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12635_ = b[535:528];
      107'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12635_ = b[543:536];
      107'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12635_ = b[551:544];
      107'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12635_ = b[559:552];
      107'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12635_ = b[567:560];
      107'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12635_ = b[575:568];
      107'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12635_ = b[583:576];
      107'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12635_ = b[591:584];
      107'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12635_ = b[599:592];
      107'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12635_ = b[607:600];
      107'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[615:608];
      107'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[623:616];
      107'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[631:624];
      107'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[639:632];
      107'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[647:640];
      107'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[655:648];
      107'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[663:656];
      107'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[671:664];
      107'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[679:672];
      107'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[687:680];
      107'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[695:688];
      107'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[703:696];
      107'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[711:704];
      107'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[719:712];
      107'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[727:720];
      107'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[735:728];
      107'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[743:736];
      107'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[751:744];
      107'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[759:752];
      107'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[767:760];
      107'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[775:768];
      107'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[783:776];
      107'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[791:784];
      107'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[799:792];
      107'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[807:800];
      107'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[815:808];
      107'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[823:816];
      107'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[831:824];
      107'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[839:832];
      107'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[847:840];
      107'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12635_ = b[855:848];
      default:
        _12635_ = a;
    endcase
  endfunction
  assign vec_data_106 = _12635_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840], data_d1[855:848] }, { _03330_, _03329_, _03328_, _03327_, _03326_, _03325_, _03324_, _03323_, _03322_, _03321_, _03320_, _03319_, _03318_, _03317_, _03316_, _03315_, _03314_, _03313_, _03312_, _03311_, _03310_, _03309_, _03308_, _03307_, _03306_, _03305_, _03304_, _03303_, _03302_, _03301_, _03300_, _03299_, _03298_, _03297_, _03296_, _03295_, _03294_, _03293_, _03292_, _03291_, _03290_, _03289_, _03288_, _03287_, _03286_, _03285_, _03284_, _03283_, _03282_, _03281_, _03280_, _03279_, _03278_, _03277_, _03276_, _03275_, _03274_, _03273_, _03272_, _03271_, _03270_, _03269_, _03268_, _03267_, _03266_, _03265_, _03264_, _03263_, _03262_, _03261_, _03260_, _03259_, _03258_, _03257_, _03256_, _03255_, _03254_, _03253_, _03252_, _03251_, _03250_, _03249_, _03248_, _03247_, _03246_, _03245_, _03244_, _03243_, _03242_, _03241_, _03240_, _03239_, _03238_, _03237_, _03236_, _03235_, _03234_, _03233_, _03232_, _03231_, _03230_, _03229_, _03228_, _03227_, _03226_, _03225_, _03224_ });
  assign _03224_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1101011;
  assign _03225_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1101010;
  assign _03226_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1101001;
  assign _03227_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1101000;
  assign _03228_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100111;
  assign _03229_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100110;
  assign _03230_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100101;
  assign _03231_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100100;
  assign _03232_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100011;
  assign _03233_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100010;
  assign _03234_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100001;
  assign _03235_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1100000;
  assign _03236_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011111;
  assign _03237_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011110;
  assign _03238_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011101;
  assign _03239_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011100;
  assign _03240_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011011;
  assign _03241_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011010;
  assign _03242_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011001;
  assign _03243_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1011000;
  assign _03244_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010111;
  assign _03245_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010110;
  assign _03246_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010101;
  assign _03247_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010100;
  assign _03248_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010011;
  assign _03249_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010010;
  assign _03250_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010001;
  assign _03251_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1010000;
  assign _03252_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001111;
  assign _03253_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001110;
  assign _03254_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001101;
  assign _03255_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001100;
  assign _03256_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001011;
  assign _03257_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001010;
  assign _03258_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001001;
  assign _03259_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1001000;
  assign _03260_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000111;
  assign _03261_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000110;
  assign _03262_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000101;
  assign _03263_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000100;
  assign _03264_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000011;
  assign _03265_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000010;
  assign _03266_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000001;
  assign _03267_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 7'b1000000;
  assign _03268_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111111;
  assign _03269_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111110;
  assign _03270_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111101;
  assign _03271_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111100;
  assign _03272_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111011;
  assign _03273_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111010;
  assign _03274_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111001;
  assign _03275_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b111000;
  assign _03276_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110111;
  assign _03277_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110110;
  assign _03278_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110101;
  assign _03279_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110100;
  assign _03280_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110011;
  assign _03281_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110010;
  assign _03282_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110001;
  assign _03283_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b110000;
  assign _03284_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101111;
  assign _03285_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101110;
  assign _03286_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101101;
  assign _03287_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101100;
  assign _03288_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101011;
  assign _03289_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101010;
  assign _03290_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101001;
  assign _03291_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b101000;
  assign _03292_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100111;
  assign _03293_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100110;
  assign _03294_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100101;
  assign _03295_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100100;
  assign _03296_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100011;
  assign _03297_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100010;
  assign _03298_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100001;
  assign _03299_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 6'b100000;
  assign _03300_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11111;
  assign _03301_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11110;
  assign _03302_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11101;
  assign _03303_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11100;
  assign _03304_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11011;
  assign _03305_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11010;
  assign _03306_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11001;
  assign _03307_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b11000;
  assign _03308_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10111;
  assign _03309_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10110;
  assign _03310_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10101;
  assign _03311_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10100;
  assign _03312_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10011;
  assign _03313_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10010;
  assign _03314_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10001;
  assign _03315_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 5'b10000;
  assign _03316_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1111;
  assign _03317_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1110;
  assign _03318_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1101;
  assign _03319_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1100;
  assign _03320_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1011;
  assign _03321_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1010;
  assign _03322_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1001;
  assign _03323_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 4'b1000;
  assign _03324_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 3'b111;
  assign _03325_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 3'b110;
  assign _03326_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 3'b101;
  assign _03327_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 3'b100;
  assign _03328_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 2'b11;
  assign _03329_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 2'b10;
  assign _03330_ = vec_sum_106_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10410" *) 1'b1;
  function [7:0] _12743_;
    input [7:0] a;
    input [847:0] b;
    input [105:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *)
    (* parallel_case *)
    casez (s)
      106'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12743_ = b[7:0];
      106'b????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12743_ = b[15:8];
      106'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12743_ = b[23:16];
      106'b??????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12743_ = b[31:24];
      106'b?????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12743_ = b[39:32];
      106'b????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12743_ = b[47:40];
      106'b???????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12743_ = b[55:48];
      106'b??????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12743_ = b[63:56];
      106'b?????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12743_ = b[71:64];
      106'b????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12743_ = b[79:72];
      106'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12743_ = b[87:80];
      106'b??????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12743_ = b[95:88];
      106'b?????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12743_ = b[103:96];
      106'b????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12743_ = b[111:104];
      106'b???????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12743_ = b[119:112];
      106'b??????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12743_ = b[127:120];
      106'b?????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12743_ = b[135:128];
      106'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12743_ = b[143:136];
      106'b???????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12743_ = b[151:144];
      106'b??????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12743_ = b[159:152];
      106'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12743_ = b[167:160];
      106'b????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12743_ = b[175:168];
      106'b???????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12743_ = b[183:176];
      106'b??????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12743_ = b[191:184];
      106'b?????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12743_ = b[199:192];
      106'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12743_ = b[207:200];
      106'b???????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12743_ = b[215:208];
      106'b??????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12743_ = b[223:216];
      106'b?????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12743_ = b[231:224];
      106'b????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12743_ = b[239:232];
      106'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12743_ = b[247:240];
      106'b??????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12743_ = b[255:248];
      106'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12743_ = b[263:256];
      106'b????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12743_ = b[271:264];
      106'b???????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12743_ = b[279:272];
      106'b??????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12743_ = b[287:280];
      106'b?????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12743_ = b[295:288];
      106'b????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12743_ = b[303:296];
      106'b???????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12743_ = b[311:304];
      106'b??????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12743_ = b[319:312];
      106'b?????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12743_ = b[327:320];
      106'b????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12743_ = b[335:328];
      106'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12743_ = b[343:336];
      106'b??????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12743_ = b[351:344];
      106'b?????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12743_ = b[359:352];
      106'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12743_ = b[367:360];
      106'b???????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12743_ = b[375:368];
      106'b??????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12743_ = b[383:376];
      106'b?????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12743_ = b[391:384];
      106'b????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12743_ = b[399:392];
      106'b???????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12743_ = b[407:400];
      106'b??????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12743_ = b[415:408];
      106'b?????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12743_ = b[423:416];
      106'b????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12743_ = b[431:424];
      106'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12743_ = b[439:432];
      106'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12743_ = b[447:440];
      106'b?????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12743_ = b[455:448];
      106'b????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12743_ = b[463:456];
      106'b???????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12743_ = b[471:464];
      106'b??????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12743_ = b[479:472];
      106'b?????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12743_ = b[487:480];
      106'b????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12743_ = b[495:488];
      106'b???????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12743_ = b[503:496];
      106'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12743_ = b[511:504];
      106'b?????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12743_ = b[519:512];
      106'b????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12743_ = b[527:520];
      106'b???????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12743_ = b[535:528];
      106'b??????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12743_ = b[543:536];
      106'b?????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12743_ = b[551:544];
      106'b????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12743_ = b[559:552];
      106'b???????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12743_ = b[567:560];
      106'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12743_ = b[575:568];
      106'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12743_ = b[583:576];
      106'b????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12743_ = b[591:584];
      106'b???????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12743_ = b[599:592];
      106'b??????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12743_ = b[607:600];
      106'b?????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[615:608];
      106'b????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[623:616];
      106'b???????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[631:624];
      106'b??????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[639:632];
      106'b?????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[647:640];
      106'b????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[655:648];
      106'b???????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[663:656];
      106'b??????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[671:664];
      106'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[679:672];
      106'b????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[687:680];
      106'b???????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[695:688];
      106'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[703:696];
      106'b?????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[711:704];
      106'b????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[719:712];
      106'b???????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[727:720];
      106'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[735:728];
      106'b?????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[743:736];
      106'b????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[751:744];
      106'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[759:752];
      106'b??????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[767:760];
      106'b?????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[775:768];
      106'b????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[783:776];
      106'b???????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[791:784];
      106'b??????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[799:792];
      106'b?????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[807:800];
      106'b????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[815:808];
      106'b???1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[823:816];
      106'b??1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[831:824];
      106'b?1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[839:832];
      106'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12743_ = b[847:840];
      default:
        _12743_ = a;
    endcase
  endfunction
  assign vec_data_105 = _12743_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832], data_d1[847:840] }, { _03436_, _03435_, _03434_, _03433_, _03432_, _03431_, _03430_, _03429_, _03428_, _03427_, _03426_, _03425_, _03424_, _03423_, _03422_, _03421_, _03420_, _03419_, _03418_, _03417_, _03416_, _03415_, _03414_, _03413_, _03412_, _03411_, _03410_, _03409_, _03408_, _03407_, _03406_, _03405_, _03404_, _03403_, _03402_, _03401_, _03400_, _03399_, _03398_, _03397_, _03396_, _03395_, _03394_, _03393_, _03392_, _03391_, _03390_, _03389_, _03388_, _03387_, _03386_, _03385_, _03384_, _03383_, _03382_, _03381_, _03380_, _03379_, _03378_, _03377_, _03376_, _03375_, _03374_, _03373_, _03372_, _03371_, _03370_, _03369_, _03368_, _03367_, _03366_, _03365_, _03364_, _03363_, _03362_, _03361_, _03360_, _03359_, _03358_, _03357_, _03356_, _03355_, _03354_, _03353_, _03352_, _03351_, _03350_, _03349_, _03348_, _03347_, _03346_, _03345_, _03344_, _03343_, _03342_, _03341_, _03340_, _03339_, _03338_, _03337_, _03336_, _03335_, _03334_, _03333_, _03332_, _03331_ });
  assign _03331_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1101010;
  assign _03332_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1101001;
  assign _03333_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1101000;
  assign _03334_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100111;
  assign _03335_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100110;
  assign _03336_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100101;
  assign _03337_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100100;
  assign _03338_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100011;
  assign _03339_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100010;
  assign _03340_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100001;
  assign _03341_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1100000;
  assign _03342_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011111;
  assign _03343_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011110;
  assign _03344_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011101;
  assign _03345_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011100;
  assign _03346_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011011;
  assign _03347_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011010;
  assign _03348_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011001;
  assign _03349_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1011000;
  assign _03350_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010111;
  assign _03351_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010110;
  assign _03352_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010101;
  assign _03353_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010100;
  assign _03354_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010011;
  assign _03355_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010010;
  assign _03356_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010001;
  assign _03357_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1010000;
  assign _03358_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001111;
  assign _03359_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001110;
  assign _03360_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001101;
  assign _03361_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001100;
  assign _03362_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001011;
  assign _03363_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001010;
  assign _03364_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001001;
  assign _03365_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1001000;
  assign _03366_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000111;
  assign _03367_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000110;
  assign _03368_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000101;
  assign _03369_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000100;
  assign _03370_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000011;
  assign _03371_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000010;
  assign _03372_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000001;
  assign _03373_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 7'b1000000;
  assign _03374_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111111;
  assign _03375_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111110;
  assign _03376_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111101;
  assign _03377_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111100;
  assign _03378_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111011;
  assign _03379_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111010;
  assign _03380_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111001;
  assign _03381_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b111000;
  assign _03382_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110111;
  assign _03383_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110110;
  assign _03384_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110101;
  assign _03385_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110100;
  assign _03386_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110011;
  assign _03387_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110010;
  assign _03388_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110001;
  assign _03389_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b110000;
  assign _03390_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101111;
  assign _03391_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101110;
  assign _03392_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101101;
  assign _03393_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101100;
  assign _03394_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101011;
  assign _03395_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101010;
  assign _03396_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101001;
  assign _03397_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b101000;
  assign _03398_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100111;
  assign _03399_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100110;
  assign _03400_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100101;
  assign _03401_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100100;
  assign _03402_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100011;
  assign _03403_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100010;
  assign _03404_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100001;
  assign _03405_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 6'b100000;
  assign _03406_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11111;
  assign _03407_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11110;
  assign _03408_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11101;
  assign _03409_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11100;
  assign _03410_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11011;
  assign _03411_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11010;
  assign _03412_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11001;
  assign _03413_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b11000;
  assign _03414_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10111;
  assign _03415_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10110;
  assign _03416_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10101;
  assign _03417_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10100;
  assign _03418_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10011;
  assign _03419_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10010;
  assign _03420_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10001;
  assign _03421_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 5'b10000;
  assign _03422_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1111;
  assign _03423_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1110;
  assign _03424_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1101;
  assign _03425_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1100;
  assign _03426_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1011;
  assign _03427_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1010;
  assign _03428_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1001;
  assign _03429_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 4'b1000;
  assign _03430_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 3'b111;
  assign _03431_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 3'b110;
  assign _03432_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 3'b101;
  assign _03433_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 3'b100;
  assign _03434_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 2'b11;
  assign _03435_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 2'b10;
  assign _03436_ = vec_sum_105_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10296" *) 1'b1;
  function [7:0] _12850_;
    input [7:0] a;
    input [839:0] b;
    input [104:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *)
    (* parallel_case *)
    casez (s)
      105'b????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12850_ = b[7:0];
      105'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12850_ = b[15:8];
      105'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12850_ = b[23:16];
      105'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12850_ = b[31:24];
      105'b????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12850_ = b[39:32];
      105'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12850_ = b[47:40];
      105'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12850_ = b[55:48];
      105'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12850_ = b[63:56];
      105'b????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12850_ = b[71:64];
      105'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12850_ = b[79:72];
      105'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12850_ = b[87:80];
      105'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12850_ = b[95:88];
      105'b????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12850_ = b[103:96];
      105'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12850_ = b[111:104];
      105'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12850_ = b[119:112];
      105'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12850_ = b[127:120];
      105'b????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12850_ = b[135:128];
      105'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12850_ = b[143:136];
      105'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12850_ = b[151:144];
      105'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12850_ = b[159:152];
      105'b????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12850_ = b[167:160];
      105'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12850_ = b[175:168];
      105'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12850_ = b[183:176];
      105'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12850_ = b[191:184];
      105'b????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12850_ = b[199:192];
      105'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12850_ = b[207:200];
      105'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12850_ = b[215:208];
      105'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12850_ = b[223:216];
      105'b????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12850_ = b[231:224];
      105'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12850_ = b[239:232];
      105'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12850_ = b[247:240];
      105'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12850_ = b[255:248];
      105'b????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12850_ = b[263:256];
      105'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12850_ = b[271:264];
      105'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12850_ = b[279:272];
      105'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12850_ = b[287:280];
      105'b????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12850_ = b[295:288];
      105'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12850_ = b[303:296];
      105'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12850_ = b[311:304];
      105'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12850_ = b[319:312];
      105'b????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12850_ = b[327:320];
      105'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12850_ = b[335:328];
      105'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12850_ = b[343:336];
      105'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12850_ = b[351:344];
      105'b????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12850_ = b[359:352];
      105'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12850_ = b[367:360];
      105'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12850_ = b[375:368];
      105'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12850_ = b[383:376];
      105'b????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12850_ = b[391:384];
      105'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12850_ = b[399:392];
      105'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12850_ = b[407:400];
      105'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12850_ = b[415:408];
      105'b????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12850_ = b[423:416];
      105'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12850_ = b[431:424];
      105'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12850_ = b[439:432];
      105'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12850_ = b[447:440];
      105'b????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12850_ = b[455:448];
      105'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12850_ = b[463:456];
      105'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12850_ = b[471:464];
      105'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12850_ = b[479:472];
      105'b????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12850_ = b[487:480];
      105'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12850_ = b[495:488];
      105'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12850_ = b[503:496];
      105'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12850_ = b[511:504];
      105'b????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12850_ = b[519:512];
      105'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12850_ = b[527:520];
      105'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12850_ = b[535:528];
      105'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12850_ = b[543:536];
      105'b????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12850_ = b[551:544];
      105'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12850_ = b[559:552];
      105'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12850_ = b[567:560];
      105'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12850_ = b[575:568];
      105'b????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12850_ = b[583:576];
      105'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12850_ = b[591:584];
      105'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12850_ = b[599:592];
      105'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12850_ = b[607:600];
      105'b????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[615:608];
      105'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[623:616];
      105'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[631:624];
      105'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[639:632];
      105'b????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[647:640];
      105'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[655:648];
      105'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[663:656];
      105'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[671:664];
      105'b????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[679:672];
      105'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[687:680];
      105'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[695:688];
      105'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[703:696];
      105'b????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[711:704];
      105'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[719:712];
      105'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[727:720];
      105'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[735:728];
      105'b????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[743:736];
      105'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[751:744];
      105'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[759:752];
      105'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[767:760];
      105'b????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[775:768];
      105'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[783:776];
      105'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[791:784];
      105'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[799:792];
      105'b????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[807:800];
      105'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[815:808];
      105'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[823:816];
      105'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[831:824];
      105'b1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12850_ = b[839:832];
      default:
        _12850_ = a;
    endcase
  endfunction
  assign vec_data_104 = _12850_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824], data_d1[839:832] }, { _03541_, _03540_, _03539_, _03538_, _03537_, _03536_, _03535_, _03534_, _03533_, _03532_, _03531_, _03530_, _03529_, _03528_, _03527_, _03526_, _03525_, _03524_, _03523_, _03522_, _03521_, _03520_, _03519_, _03518_, _03517_, _03516_, _03515_, _03514_, _03513_, _03512_, _03511_, _03510_, _03509_, _03508_, _03507_, _03506_, _03505_, _03504_, _03503_, _03502_, _03501_, _03500_, _03499_, _03498_, _03497_, _03496_, _03495_, _03494_, _03493_, _03492_, _03491_, _03490_, _03489_, _03488_, _03487_, _03486_, _03485_, _03484_, _03483_, _03482_, _03481_, _03480_, _03479_, _03478_, _03477_, _03476_, _03475_, _03474_, _03473_, _03472_, _03471_, _03470_, _03469_, _03468_, _03467_, _03466_, _03465_, _03464_, _03463_, _03462_, _03461_, _03460_, _03459_, _03458_, _03457_, _03456_, _03455_, _03454_, _03453_, _03452_, _03451_, _03450_, _03449_, _03448_, _03447_, _03446_, _03445_, _03444_, _03443_, _03442_, _03441_, _03440_, _03439_, _03438_, _03437_ });
  assign _03437_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1101001;
  assign _03438_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1101000;
  assign _03439_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100111;
  assign _03440_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100110;
  assign _03441_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100101;
  assign _03442_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100100;
  assign _03443_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100011;
  assign _03444_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100010;
  assign _03445_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100001;
  assign _03446_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1100000;
  assign _03447_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011111;
  assign _03448_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011110;
  assign _03449_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011101;
  assign _03450_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011100;
  assign _03451_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011011;
  assign _03452_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011010;
  assign _03453_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011001;
  assign _03454_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1011000;
  assign _03455_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010111;
  assign _03456_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010110;
  assign _03457_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010101;
  assign _03458_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010100;
  assign _03459_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010011;
  assign _03460_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010010;
  assign _03461_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010001;
  assign _03462_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1010000;
  assign _03463_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001111;
  assign _03464_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001110;
  assign _03465_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001101;
  assign _03466_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001100;
  assign _03467_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001011;
  assign _03468_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001010;
  assign _03469_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001001;
  assign _03470_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1001000;
  assign _03471_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000111;
  assign _03472_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000110;
  assign _03473_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000101;
  assign _03474_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000100;
  assign _03475_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000011;
  assign _03476_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000010;
  assign _03477_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000001;
  assign _03478_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 7'b1000000;
  assign _03479_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111111;
  assign _03480_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111110;
  assign _03481_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111101;
  assign _03482_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111100;
  assign _03483_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111011;
  assign _03484_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111010;
  assign _03485_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111001;
  assign _03486_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b111000;
  assign _03487_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110111;
  assign _03488_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110110;
  assign _03489_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110101;
  assign _03490_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110100;
  assign _03491_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110011;
  assign _03492_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10233|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110010;
  assign _03493_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110001;
  assign _03494_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b110000;
  assign _03495_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101111;
  assign _03496_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101110;
  assign _03497_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101101;
  assign _03498_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101100;
  assign _03499_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101011;
  assign _03500_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101010;
  assign _03501_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101001;
  assign _03502_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b101000;
  assign _03503_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100111;
  assign _03504_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100110;
  assign _03505_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100101;
  assign _03506_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100100;
  assign _03507_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100011;
  assign _03508_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100010;
  assign _03509_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100001;
  assign _03510_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 6'b100000;
  assign _03511_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11111;
  assign _03512_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11110;
  assign _03513_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11101;
  assign _03514_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11100;
  assign _03515_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11011;
  assign _03516_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11010;
  assign _03517_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11001;
  assign _03518_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b11000;
  assign _03519_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10111;
  assign _03520_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10110;
  assign _03521_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10101;
  assign _03522_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10100;
  assign _03523_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10011;
  assign _03524_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10010;
  assign _03525_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10001;
  assign _03526_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 5'b10000;
  assign _03527_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1111;
  assign _03528_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1110;
  assign _03529_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1101;
  assign _03530_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1100;
  assign _03531_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1011;
  assign _03532_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1010;
  assign _03533_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1001;
  assign _03534_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 4'b1000;
  assign _03535_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 3'b111;
  assign _03536_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 3'b110;
  assign _03537_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 3'b101;
  assign _03538_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 3'b100;
  assign _03539_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 2'b11;
  assign _03540_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 2'b10;
  assign _03541_ = vec_sum_104_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10183" *) 1'b1;
  function [7:0] _12956_;
    input [7:0] a;
    input [831:0] b;
    input [103:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *)
    (* parallel_case *)
    casez (s)
      104'b???????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _12956_ = b[7:0];
      104'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _12956_ = b[15:8];
      104'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _12956_ = b[23:16];
      104'b????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _12956_ = b[31:24];
      104'b???????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _12956_ = b[39:32];
      104'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _12956_ = b[47:40];
      104'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _12956_ = b[55:48];
      104'b????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _12956_ = b[63:56];
      104'b???????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _12956_ = b[71:64];
      104'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _12956_ = b[79:72];
      104'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _12956_ = b[87:80];
      104'b????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _12956_ = b[95:88];
      104'b???????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _12956_ = b[103:96];
      104'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _12956_ = b[111:104];
      104'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _12956_ = b[119:112];
      104'b????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _12956_ = b[127:120];
      104'b???????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _12956_ = b[135:128];
      104'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _12956_ = b[143:136];
      104'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _12956_ = b[151:144];
      104'b????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _12956_ = b[159:152];
      104'b???????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _12956_ = b[167:160];
      104'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _12956_ = b[175:168];
      104'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _12956_ = b[183:176];
      104'b????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _12956_ = b[191:184];
      104'b???????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _12956_ = b[199:192];
      104'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _12956_ = b[207:200];
      104'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _12956_ = b[215:208];
      104'b????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _12956_ = b[223:216];
      104'b???????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _12956_ = b[231:224];
      104'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _12956_ = b[239:232];
      104'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _12956_ = b[247:240];
      104'b????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _12956_ = b[255:248];
      104'b???????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _12956_ = b[263:256];
      104'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _12956_ = b[271:264];
      104'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _12956_ = b[279:272];
      104'b????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _12956_ = b[287:280];
      104'b???????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _12956_ = b[295:288];
      104'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _12956_ = b[303:296];
      104'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _12956_ = b[311:304];
      104'b????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _12956_ = b[319:312];
      104'b???????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _12956_ = b[327:320];
      104'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _12956_ = b[335:328];
      104'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _12956_ = b[343:336];
      104'b????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _12956_ = b[351:344];
      104'b???????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _12956_ = b[359:352];
      104'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _12956_ = b[367:360];
      104'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _12956_ = b[375:368];
      104'b????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _12956_ = b[383:376];
      104'b???????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _12956_ = b[391:384];
      104'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _12956_ = b[399:392];
      104'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _12956_ = b[407:400];
      104'b????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _12956_ = b[415:408];
      104'b???????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _12956_ = b[423:416];
      104'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _12956_ = b[431:424];
      104'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _12956_ = b[439:432];
      104'b????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _12956_ = b[447:440];
      104'b???????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _12956_ = b[455:448];
      104'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _12956_ = b[463:456];
      104'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _12956_ = b[471:464];
      104'b????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _12956_ = b[479:472];
      104'b???????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _12956_ = b[487:480];
      104'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _12956_ = b[495:488];
      104'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _12956_ = b[503:496];
      104'b????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _12956_ = b[511:504];
      104'b???????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _12956_ = b[519:512];
      104'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _12956_ = b[527:520];
      104'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _12956_ = b[535:528];
      104'b????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _12956_ = b[543:536];
      104'b???????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _12956_ = b[551:544];
      104'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _12956_ = b[559:552];
      104'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _12956_ = b[567:560];
      104'b????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _12956_ = b[575:568];
      104'b???????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _12956_ = b[583:576];
      104'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _12956_ = b[591:584];
      104'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _12956_ = b[599:592];
      104'b????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _12956_ = b[607:600];
      104'b???????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[615:608];
      104'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[623:616];
      104'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[631:624];
      104'b????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[639:632];
      104'b???????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[647:640];
      104'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[655:648];
      104'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[663:656];
      104'b????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[671:664];
      104'b???????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[679:672];
      104'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[687:680];
      104'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[695:688];
      104'b????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[703:696];
      104'b???????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[711:704];
      104'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[719:712];
      104'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[727:720];
      104'b????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[735:728];
      104'b???????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[743:736];
      104'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[751:744];
      104'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[759:752];
      104'b????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[767:760];
      104'b???????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[775:768];
      104'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[783:776];
      104'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[791:784];
      104'b????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[799:792];
      104'b???1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[807:800];
      104'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[815:808];
      104'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[823:816];
      104'b1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _12956_ = b[831:824];
      default:
        _12956_ = a;
    endcase
  endfunction
  assign vec_data_103 = _12956_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816], data_d1[831:824] }, { _03645_, _03644_, _03643_, _03642_, _03641_, _03640_, _03639_, _03638_, _03637_, _03636_, _03635_, _03634_, _03633_, _03632_, _03631_, _03630_, _03629_, _03628_, _03627_, _03626_, _03625_, _03624_, _03623_, _03622_, _03621_, _03620_, _03619_, _03618_, _03617_, _03616_, _03615_, _03614_, _03613_, _03612_, _03611_, _03610_, _03609_, _03608_, _03607_, _03606_, _03605_, _03604_, _03603_, _03602_, _03601_, _03600_, _03599_, _03598_, _03597_, _03596_, _03595_, _03594_, _03593_, _03592_, _03591_, _03590_, _03589_, _03588_, _03587_, _03586_, _03585_, _03584_, _03583_, _03582_, _03581_, _03580_, _03579_, _03578_, _03577_, _03576_, _03575_, _03574_, _03573_, _03572_, _03571_, _03570_, _03569_, _03568_, _03567_, _03566_, _03565_, _03564_, _03563_, _03562_, _03561_, _03560_, _03559_, _03558_, _03557_, _03556_, _03555_, _03554_, _03553_, _03552_, _03551_, _03550_, _03549_, _03548_, _03547_, _03546_, _03545_, _03544_, _03543_, _03542_ });
  assign _03542_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1101000;
  assign _03543_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100111;
  assign _03544_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100110;
  assign _03545_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100101;
  assign _03546_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100100;
  assign _03547_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100011;
  assign _03548_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100010;
  assign _03549_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100001;
  assign _03550_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1100000;
  assign _03551_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011111;
  assign _03552_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011110;
  assign _03553_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011101;
  assign _03554_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011100;
  assign _03555_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011011;
  assign _03556_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011010;
  assign _03557_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011001;
  assign _03558_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1011000;
  assign _03559_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010111;
  assign _03560_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010110;
  assign _03561_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010101;
  assign _03562_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010100;
  assign _03563_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010011;
  assign _03564_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010010;
  assign _03565_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010001;
  assign _03566_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1010000;
  assign _03567_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001111;
  assign _03568_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001110;
  assign _03569_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001101;
  assign _03570_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001100;
  assign _03571_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001011;
  assign _03572_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001010;
  assign _03573_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001001;
  assign _03574_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1001000;
  assign _03575_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000111;
  assign _03576_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000110;
  assign _03577_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000101;
  assign _03578_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000100;
  assign _03579_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000011;
  assign _03580_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000010;
  assign _03581_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000001;
  assign _03582_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 7'b1000000;
  assign _03583_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111111;
  assign _03584_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111110;
  assign _03585_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111101;
  assign _03586_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111100;
  assign _03587_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111011;
  assign _03588_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111010;
  assign _03589_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111001;
  assign _03590_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b111000;
  assign _03591_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110111;
  assign _03592_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110110;
  assign _03593_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110101;
  assign _03594_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110100;
  assign _03595_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110011;
  assign _03596_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110010;
  assign _03597_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110001;
  assign _03598_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b110000;
  assign _03599_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101111;
  assign _03600_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101110;
  assign _03601_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101101;
  assign _03602_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101100;
  assign _03603_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101011;
  assign _03604_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101010;
  assign _03605_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101001;
  assign _03606_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b101000;
  assign _03607_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100111;
  assign _03608_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100110;
  assign _03609_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100101;
  assign _03610_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100100;
  assign _03611_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100011;
  assign _03612_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100010;
  assign _03613_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100001;
  assign _03614_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 6'b100000;
  assign _03615_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11111;
  assign _03616_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11110;
  assign _03617_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11101;
  assign _03618_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11100;
  assign _03619_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11011;
  assign _03620_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11010;
  assign _03621_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11001;
  assign _03622_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b11000;
  assign _03623_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10111;
  assign _03624_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10110;
  assign _03625_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10101;
  assign _03626_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10100;
  assign _03627_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10011;
  assign _03628_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10010;
  assign _03629_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10001;
  assign _03630_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 5'b10000;
  assign _03631_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1111;
  assign _03632_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1110;
  assign _03633_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1101;
  assign _03634_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1100;
  assign _03635_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1011;
  assign _03636_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1010;
  assign _03637_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1001;
  assign _03638_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 4'b1000;
  assign _03639_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 3'b111;
  assign _03640_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 3'b110;
  assign _03641_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 3'b101;
  assign _03642_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 3'b100;
  assign _03643_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 2'b11;
  assign _03644_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 2'b10;
  assign _03645_ = vec_sum_103_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10071" *) 1'b1;
  function [7:0] _13061_;
    input [7:0] a;
    input [823:0] b;
    input [102:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *)
    (* parallel_case *)
    casez (s)
      103'b??????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13061_ = b[7:0];
      103'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13061_ = b[15:8];
      103'b????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13061_ = b[23:16];
      103'b???????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13061_ = b[31:24];
      103'b??????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13061_ = b[39:32];
      103'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13061_ = b[47:40];
      103'b????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13061_ = b[55:48];
      103'b???????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13061_ = b[63:56];
      103'b??????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13061_ = b[71:64];
      103'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13061_ = b[79:72];
      103'b????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13061_ = b[87:80];
      103'b???????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13061_ = b[95:88];
      103'b??????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13061_ = b[103:96];
      103'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13061_ = b[111:104];
      103'b????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13061_ = b[119:112];
      103'b???????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13061_ = b[127:120];
      103'b??????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13061_ = b[135:128];
      103'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13061_ = b[143:136];
      103'b????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13061_ = b[151:144];
      103'b???????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13061_ = b[159:152];
      103'b??????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13061_ = b[167:160];
      103'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13061_ = b[175:168];
      103'b????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13061_ = b[183:176];
      103'b???????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13061_ = b[191:184];
      103'b??????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13061_ = b[199:192];
      103'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13061_ = b[207:200];
      103'b????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13061_ = b[215:208];
      103'b???????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13061_ = b[223:216];
      103'b??????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13061_ = b[231:224];
      103'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13061_ = b[239:232];
      103'b????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13061_ = b[247:240];
      103'b???????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13061_ = b[255:248];
      103'b??????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13061_ = b[263:256];
      103'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13061_ = b[271:264];
      103'b????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13061_ = b[279:272];
      103'b???????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13061_ = b[287:280];
      103'b??????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13061_ = b[295:288];
      103'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13061_ = b[303:296];
      103'b????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13061_ = b[311:304];
      103'b???????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13061_ = b[319:312];
      103'b??????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13061_ = b[327:320];
      103'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13061_ = b[335:328];
      103'b????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13061_ = b[343:336];
      103'b???????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13061_ = b[351:344];
      103'b??????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13061_ = b[359:352];
      103'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13061_ = b[367:360];
      103'b????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13061_ = b[375:368];
      103'b???????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13061_ = b[383:376];
      103'b??????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13061_ = b[391:384];
      103'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13061_ = b[399:392];
      103'b????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13061_ = b[407:400];
      103'b???????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13061_ = b[415:408];
      103'b??????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13061_ = b[423:416];
      103'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13061_ = b[431:424];
      103'b????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13061_ = b[439:432];
      103'b???????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13061_ = b[447:440];
      103'b??????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13061_ = b[455:448];
      103'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13061_ = b[463:456];
      103'b????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13061_ = b[471:464];
      103'b???????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13061_ = b[479:472];
      103'b??????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13061_ = b[487:480];
      103'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13061_ = b[495:488];
      103'b????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13061_ = b[503:496];
      103'b???????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13061_ = b[511:504];
      103'b??????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13061_ = b[519:512];
      103'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13061_ = b[527:520];
      103'b????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13061_ = b[535:528];
      103'b???????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13061_ = b[543:536];
      103'b??????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13061_ = b[551:544];
      103'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13061_ = b[559:552];
      103'b????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13061_ = b[567:560];
      103'b???????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13061_ = b[575:568];
      103'b??????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13061_ = b[583:576];
      103'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13061_ = b[591:584];
      103'b????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13061_ = b[599:592];
      103'b???????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13061_ = b[607:600];
      103'b??????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[615:608];
      103'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[623:616];
      103'b????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[631:624];
      103'b???????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[639:632];
      103'b??????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[647:640];
      103'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[655:648];
      103'b????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[663:656];
      103'b???????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[671:664];
      103'b??????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[679:672];
      103'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[687:680];
      103'b????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[695:688];
      103'b???????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[703:696];
      103'b??????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[711:704];
      103'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[719:712];
      103'b????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[727:720];
      103'b???????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[735:728];
      103'b??????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[743:736];
      103'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[751:744];
      103'b????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[759:752];
      103'b???????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[767:760];
      103'b??????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[775:768];
      103'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[783:776];
      103'b????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[791:784];
      103'b???1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[799:792];
      103'b??1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[807:800];
      103'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[815:808];
      103'b1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13061_ = b[823:816];
      default:
        _13061_ = a;
    endcase
  endfunction
  assign vec_data_102 = _13061_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808], data_d1[823:816] }, { _03748_, _03747_, _03746_, _03745_, _03744_, _03743_, _03742_, _03741_, _03740_, _03739_, _03738_, _03737_, _03736_, _03735_, _03734_, _03733_, _03732_, _03731_, _03730_, _03729_, _03728_, _03727_, _03726_, _03725_, _03724_, _03723_, _03722_, _03721_, _03720_, _03719_, _03718_, _03717_, _03716_, _03715_, _03714_, _03713_, _03712_, _03711_, _03710_, _03709_, _03708_, _03707_, _03706_, _03705_, _03704_, _03703_, _03702_, _03701_, _03700_, _03699_, _03698_, _03697_, _03696_, _03695_, _03694_, _03693_, _03692_, _03691_, _03690_, _03689_, _03688_, _03687_, _03686_, _03685_, _03684_, _03683_, _03682_, _03681_, _03680_, _03679_, _03678_, _03677_, _03676_, _03675_, _03674_, _03673_, _03672_, _03671_, _03670_, _03669_, _03668_, _03667_, _03666_, _03665_, _03664_, _03663_, _03662_, _03661_, _03660_, _03659_, _03658_, _03657_, _03656_, _03655_, _03654_, _03653_, _03652_, _03651_, _03650_, _03649_, _03648_, _03647_, _03646_ });
  assign _03646_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100111;
  assign _03647_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100110;
  assign _03648_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100101;
  assign _03649_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100100;
  assign _03650_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100011;
  assign _03651_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100010;
  assign _03652_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100001;
  assign _03653_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1100000;
  assign _03654_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011111;
  assign _03655_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011110;
  assign _03656_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011101;
  assign _03657_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011100;
  assign _03658_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011011;
  assign _03659_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011010;
  assign _03660_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011001;
  assign _03661_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1011000;
  assign _03662_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010111;
  assign _03663_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010110;
  assign _03664_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010101;
  assign _03665_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010100;
  assign _03666_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010011;
  assign _03667_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010010;
  assign _03668_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010001;
  assign _03669_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1010000;
  assign _03670_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001111;
  assign _03671_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001110;
  assign _03672_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001101;
  assign _03673_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001100;
  assign _03674_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001011;
  assign _03675_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001010;
  assign _03676_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001001;
  assign _03677_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1001000;
  assign _03678_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000111;
  assign _03679_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000110;
  assign _03680_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000101;
  assign _03681_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000100;
  assign _03682_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000011;
  assign _03683_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000010;
  assign _03684_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000001;
  assign _03685_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 7'b1000000;
  assign _03686_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111111;
  assign _03687_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111110;
  assign _03688_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111101;
  assign _03689_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111100;
  assign _03690_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111011;
  assign _03691_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111010;
  assign _03692_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111001;
  assign _03693_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b111000;
  assign _03694_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110111;
  assign _03695_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110110;
  assign _03696_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110101;
  assign _03697_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110100;
  assign _03698_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110011;
  assign _03699_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110010;
  assign _03700_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110001;
  assign _03701_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b110000;
  assign _03702_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101111;
  assign _03703_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101110;
  assign _03704_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101101;
  assign _03705_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101100;
  assign _03706_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101011;
  assign _03707_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101010;
  assign _03708_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101001;
  assign _03709_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:10000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b101000;
  assign _03710_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100111;
  assign _03711_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100110;
  assign _03712_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100101;
  assign _03713_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100100;
  assign _03714_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100011;
  assign _03715_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100010;
  assign _03716_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100001;
  assign _03717_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 6'b100000;
  assign _03718_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11111;
  assign _03719_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11110;
  assign _03720_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11101;
  assign _03721_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11100;
  assign _03722_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11011;
  assign _03723_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11010;
  assign _03724_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11001;
  assign _03725_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b11000;
  assign _03726_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10111;
  assign _03727_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10110;
  assign _03728_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10101;
  assign _03729_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10100;
  assign _03730_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10011;
  assign _03731_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10010;
  assign _03732_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10001;
  assign _03733_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 5'b10000;
  assign _03734_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1111;
  assign _03735_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1110;
  assign _03736_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1101;
  assign _03737_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1100;
  assign _03738_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1011;
  assign _03739_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1010;
  assign _03740_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1001;
  assign _03741_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 4'b1000;
  assign _03742_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 3'b111;
  assign _03743_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 3'b110;
  assign _03744_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 3'b101;
  assign _03745_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 3'b100;
  assign _03746_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 2'b11;
  assign _03747_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 2'b10;
  assign _03748_ = vec_sum_102_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9960" *) 1'b1;
  function [7:0] _13165_;
    input [7:0] a;
    input [815:0] b;
    input [101:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *)
    (* parallel_case *)
    casez (s)
      102'b?????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13165_ = b[7:0];
      102'b????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13165_ = b[15:8];
      102'b???????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13165_ = b[23:16];
      102'b??????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13165_ = b[31:24];
      102'b?????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13165_ = b[39:32];
      102'b????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13165_ = b[47:40];
      102'b???????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13165_ = b[55:48];
      102'b??????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13165_ = b[63:56];
      102'b?????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13165_ = b[71:64];
      102'b????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13165_ = b[79:72];
      102'b???????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13165_ = b[87:80];
      102'b??????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13165_ = b[95:88];
      102'b?????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13165_ = b[103:96];
      102'b????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13165_ = b[111:104];
      102'b???????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13165_ = b[119:112];
      102'b??????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13165_ = b[127:120];
      102'b?????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13165_ = b[135:128];
      102'b????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13165_ = b[143:136];
      102'b???????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13165_ = b[151:144];
      102'b??????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13165_ = b[159:152];
      102'b?????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13165_ = b[167:160];
      102'b????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13165_ = b[175:168];
      102'b???????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13165_ = b[183:176];
      102'b??????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13165_ = b[191:184];
      102'b?????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13165_ = b[199:192];
      102'b????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13165_ = b[207:200];
      102'b???????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13165_ = b[215:208];
      102'b??????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13165_ = b[223:216];
      102'b?????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13165_ = b[231:224];
      102'b????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13165_ = b[239:232];
      102'b???????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13165_ = b[247:240];
      102'b??????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13165_ = b[255:248];
      102'b?????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13165_ = b[263:256];
      102'b????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13165_ = b[271:264];
      102'b???????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13165_ = b[279:272];
      102'b??????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13165_ = b[287:280];
      102'b?????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13165_ = b[295:288];
      102'b????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13165_ = b[303:296];
      102'b???????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13165_ = b[311:304];
      102'b??????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13165_ = b[319:312];
      102'b?????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13165_ = b[327:320];
      102'b????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13165_ = b[335:328];
      102'b???????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13165_ = b[343:336];
      102'b??????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13165_ = b[351:344];
      102'b?????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13165_ = b[359:352];
      102'b????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13165_ = b[367:360];
      102'b???????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13165_ = b[375:368];
      102'b??????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13165_ = b[383:376];
      102'b?????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13165_ = b[391:384];
      102'b????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13165_ = b[399:392];
      102'b???????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13165_ = b[407:400];
      102'b??????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13165_ = b[415:408];
      102'b?????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13165_ = b[423:416];
      102'b????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13165_ = b[431:424];
      102'b???????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13165_ = b[439:432];
      102'b??????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13165_ = b[447:440];
      102'b?????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13165_ = b[455:448];
      102'b????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13165_ = b[463:456];
      102'b???????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13165_ = b[471:464];
      102'b??????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13165_ = b[479:472];
      102'b?????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13165_ = b[487:480];
      102'b????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13165_ = b[495:488];
      102'b???????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13165_ = b[503:496];
      102'b??????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13165_ = b[511:504];
      102'b?????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13165_ = b[519:512];
      102'b????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13165_ = b[527:520];
      102'b???????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13165_ = b[535:528];
      102'b??????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13165_ = b[543:536];
      102'b?????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13165_ = b[551:544];
      102'b????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13165_ = b[559:552];
      102'b???????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13165_ = b[567:560];
      102'b??????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13165_ = b[575:568];
      102'b?????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13165_ = b[583:576];
      102'b????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13165_ = b[591:584];
      102'b???????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13165_ = b[599:592];
      102'b??????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13165_ = b[607:600];
      102'b?????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[615:608];
      102'b????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[623:616];
      102'b???????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[631:624];
      102'b??????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[639:632];
      102'b?????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[647:640];
      102'b????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[655:648];
      102'b???????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[663:656];
      102'b??????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[671:664];
      102'b?????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[679:672];
      102'b????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[687:680];
      102'b???????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[695:688];
      102'b??????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[703:696];
      102'b?????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[711:704];
      102'b????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[719:712];
      102'b???????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[727:720];
      102'b??????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[735:728];
      102'b?????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[743:736];
      102'b????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[751:744];
      102'b???????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[759:752];
      102'b??????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[767:760];
      102'b?????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[775:768];
      102'b????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[783:776];
      102'b???1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[791:784];
      102'b??1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[799:792];
      102'b?1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[807:800];
      102'b1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13165_ = b[815:808];
      default:
        _13165_ = a;
    endcase
  endfunction
  assign vec_data_101 = _13165_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800], data_d1[815:808] }, { _03850_, _03849_, _03848_, _03847_, _03846_, _03845_, _03844_, _03843_, _03842_, _03841_, _03840_, _03839_, _03838_, _03837_, _03836_, _03835_, _03834_, _03833_, _03832_, _03831_, _03830_, _03829_, _03828_, _03827_, _03826_, _03825_, _03824_, _03823_, _03822_, _03821_, _03820_, _03819_, _03818_, _03817_, _03816_, _03815_, _03814_, _03813_, _03812_, _03811_, _03810_, _03809_, _03808_, _03807_, _03806_, _03805_, _03804_, _03803_, _03802_, _03801_, _03800_, _03799_, _03798_, _03797_, _03796_, _03795_, _03794_, _03793_, _03792_, _03791_, _03790_, _03789_, _03788_, _03787_, _03786_, _03785_, _03784_, _03783_, _03782_, _03781_, _03780_, _03779_, _03778_, _03777_, _03776_, _03775_, _03774_, _03773_, _03772_, _03771_, _03770_, _03769_, _03768_, _03767_, _03766_, _03765_, _03764_, _03763_, _03762_, _03761_, _03760_, _03759_, _03758_, _03757_, _03756_, _03755_, _03754_, _03753_, _03752_, _03751_, _03750_, _03749_ });
  assign _03749_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100110;
  assign _03750_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100101;
  assign _03751_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100100;
  assign _03752_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100011;
  assign _03753_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100010;
  assign _03754_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100001;
  assign _03755_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1100000;
  assign _03756_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011111;
  assign _03757_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011110;
  assign _03758_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011101;
  assign _03759_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011100;
  assign _03760_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011011;
  assign _03761_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011010;
  assign _03762_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011001;
  assign _03763_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1011000;
  assign _03764_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010111;
  assign _03765_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010110;
  assign _03766_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010101;
  assign _03767_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010100;
  assign _03768_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010011;
  assign _03769_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010010;
  assign _03770_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010001;
  assign _03771_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1010000;
  assign _03772_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001111;
  assign _03773_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001110;
  assign _03774_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001101;
  assign _03775_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001100;
  assign _03776_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001011;
  assign _03777_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001010;
  assign _03778_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001001;
  assign _03779_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1001000;
  assign _03780_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000111;
  assign _03781_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000110;
  assign _03782_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000101;
  assign _03783_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000100;
  assign _03784_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000011;
  assign _03785_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000010;
  assign _03786_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000001;
  assign _03787_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 7'b1000000;
  assign _03788_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111111;
  assign _03789_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111110;
  assign _03790_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111101;
  assign _03791_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111100;
  assign _03792_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111011;
  assign _03793_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111010;
  assign _03794_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111001;
  assign _03795_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b111000;
  assign _03796_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110111;
  assign _03797_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110110;
  assign _03798_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110101;
  assign _03799_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110100;
  assign _03800_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110011;
  assign _03801_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110010;
  assign _03802_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110001;
  assign _03803_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b110000;
  assign _03804_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101111;
  assign _03805_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101110;
  assign _03806_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101101;
  assign _03807_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101100;
  assign _03808_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101011;
  assign _03809_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101010;
  assign _03810_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101001;
  assign _03811_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b101000;
  assign _03812_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100111;
  assign _03813_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100110;
  assign _03814_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100101;
  assign _03815_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100100;
  assign _03816_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100011;
  assign _03817_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100010;
  assign _03818_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100001;
  assign _03819_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 6'b100000;
  assign _03820_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11111;
  assign _03821_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11110;
  assign _03822_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11101;
  assign _03823_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11100;
  assign _03824_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11011;
  assign _03825_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11010;
  assign _03826_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11001;
  assign _03827_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b11000;
  assign _03828_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10111;
  assign _03829_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10110;
  assign _03830_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10101;
  assign _03831_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10100;
  assign _03832_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10011;
  assign _03833_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10010;
  assign _03834_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10001;
  assign _03835_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 5'b10000;
  assign _03836_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1111;
  assign _03837_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1110;
  assign _03838_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1101;
  assign _03839_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1100;
  assign _03840_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1011;
  assign _03841_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1010;
  assign _03842_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1001;
  assign _03843_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 4'b1000;
  assign _03844_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 3'b111;
  assign _03845_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 3'b110;
  assign _03846_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 3'b101;
  assign _03847_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 3'b100;
  assign _03848_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 2'b11;
  assign _03849_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 2'b10;
  assign _03850_ = vec_sum_101_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9850" *) 1'b1;
  function [7:0] _13268_;
    input [7:0] a;
    input [807:0] b;
    input [100:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *)
    (* parallel_case *)
    casez (s)
      101'b????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13268_ = b[7:0];
      101'b???????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13268_ = b[15:8];
      101'b??????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13268_ = b[23:16];
      101'b?????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13268_ = b[31:24];
      101'b????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13268_ = b[39:32];
      101'b???????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13268_ = b[47:40];
      101'b??????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13268_ = b[55:48];
      101'b?????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13268_ = b[63:56];
      101'b????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13268_ = b[71:64];
      101'b???????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13268_ = b[79:72];
      101'b??????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13268_ = b[87:80];
      101'b?????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13268_ = b[95:88];
      101'b????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13268_ = b[103:96];
      101'b???????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13268_ = b[111:104];
      101'b??????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13268_ = b[119:112];
      101'b?????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13268_ = b[127:120];
      101'b????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13268_ = b[135:128];
      101'b???????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13268_ = b[143:136];
      101'b??????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13268_ = b[151:144];
      101'b?????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13268_ = b[159:152];
      101'b????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13268_ = b[167:160];
      101'b???????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13268_ = b[175:168];
      101'b??????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13268_ = b[183:176];
      101'b?????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13268_ = b[191:184];
      101'b????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13268_ = b[199:192];
      101'b???????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13268_ = b[207:200];
      101'b??????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13268_ = b[215:208];
      101'b?????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13268_ = b[223:216];
      101'b????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13268_ = b[231:224];
      101'b???????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13268_ = b[239:232];
      101'b??????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13268_ = b[247:240];
      101'b?????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13268_ = b[255:248];
      101'b????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13268_ = b[263:256];
      101'b???????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13268_ = b[271:264];
      101'b??????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13268_ = b[279:272];
      101'b?????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13268_ = b[287:280];
      101'b????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13268_ = b[295:288];
      101'b???????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13268_ = b[303:296];
      101'b??????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13268_ = b[311:304];
      101'b?????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13268_ = b[319:312];
      101'b????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13268_ = b[327:320];
      101'b???????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13268_ = b[335:328];
      101'b??????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13268_ = b[343:336];
      101'b?????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13268_ = b[351:344];
      101'b????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13268_ = b[359:352];
      101'b???????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13268_ = b[367:360];
      101'b??????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13268_ = b[375:368];
      101'b?????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13268_ = b[383:376];
      101'b????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13268_ = b[391:384];
      101'b???????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13268_ = b[399:392];
      101'b??????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13268_ = b[407:400];
      101'b?????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13268_ = b[415:408];
      101'b????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13268_ = b[423:416];
      101'b???????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13268_ = b[431:424];
      101'b??????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13268_ = b[439:432];
      101'b?????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13268_ = b[447:440];
      101'b????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13268_ = b[455:448];
      101'b???????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13268_ = b[463:456];
      101'b??????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13268_ = b[471:464];
      101'b?????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13268_ = b[479:472];
      101'b????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13268_ = b[487:480];
      101'b???????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13268_ = b[495:488];
      101'b??????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13268_ = b[503:496];
      101'b?????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13268_ = b[511:504];
      101'b????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13268_ = b[519:512];
      101'b???????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13268_ = b[527:520];
      101'b??????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13268_ = b[535:528];
      101'b?????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13268_ = b[543:536];
      101'b????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13268_ = b[551:544];
      101'b???????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13268_ = b[559:552];
      101'b??????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13268_ = b[567:560];
      101'b?????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13268_ = b[575:568];
      101'b????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13268_ = b[583:576];
      101'b???????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13268_ = b[591:584];
      101'b??????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13268_ = b[599:592];
      101'b?????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13268_ = b[607:600];
      101'b????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[615:608];
      101'b???????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[623:616];
      101'b??????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[631:624];
      101'b?????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[639:632];
      101'b????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[647:640];
      101'b???????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[655:648];
      101'b??????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[663:656];
      101'b?????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[671:664];
      101'b????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[679:672];
      101'b???????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[687:680];
      101'b??????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[695:688];
      101'b?????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[703:696];
      101'b????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[711:704];
      101'b???????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[719:712];
      101'b??????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[727:720];
      101'b?????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[735:728];
      101'b????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[743:736];
      101'b???????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[751:744];
      101'b??????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[759:752];
      101'b?????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[767:760];
      101'b????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[775:768];
      101'b???1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[783:776];
      101'b??1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[791:784];
      101'b?1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[799:792];
      101'b1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _13268_ = b[807:800];
      default:
        _13268_ = a;
    endcase
  endfunction
  assign vec_data_100 = _13268_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792], data_d1[807:800] }, { _03951_, _03950_, _03949_, _03948_, _03947_, _03946_, _03945_, _03944_, _03943_, _03942_, _03941_, _03940_, _03939_, _03938_, _03937_, _03936_, _03935_, _03934_, _03933_, _03932_, _03931_, _03930_, _03929_, _03928_, _03927_, _03926_, _03925_, _03924_, _03923_, _03922_, _03921_, _03920_, _03919_, _03918_, _03917_, _03916_, _03915_, _03914_, _03913_, _03912_, _03911_, _03910_, _03909_, _03908_, _03907_, _03906_, _03905_, _03904_, _03903_, _03902_, _03901_, _03900_, _03899_, _03898_, _03897_, _03896_, _03895_, _03894_, _03893_, _03892_, _03891_, _03890_, _03889_, _03888_, _03887_, _03886_, _03885_, _03884_, _03883_, _03882_, _03881_, _03880_, _03879_, _03878_, _03877_, _03876_, _03875_, _03874_, _03873_, _03872_, _03871_, _03870_, _03869_, _03868_, _03867_, _03866_, _03865_, _03864_, _03863_, _03862_, _03861_, _03860_, _03859_, _03858_, _03857_, _03856_, _03855_, _03854_, _03853_, _03852_, _03851_ });
  assign _03851_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100101;
  assign _03852_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100100;
  assign _03853_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100011;
  assign _03854_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100010;
  assign _03855_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100001;
  assign _03856_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1100000;
  assign _03857_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011111;
  assign _03858_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011110;
  assign _03859_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011101;
  assign _03860_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011100;
  assign _03861_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011011;
  assign _03862_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011010;
  assign _03863_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011001;
  assign _03864_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1011000;
  assign _03865_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010111;
  assign _03866_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010110;
  assign _03867_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010101;
  assign _03868_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010100;
  assign _03869_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010011;
  assign _03870_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010010;
  assign _03871_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010001;
  assign _03872_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1010000;
  assign _03873_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001111;
  assign _03874_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001110;
  assign _03875_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001101;
  assign _03876_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001100;
  assign _03877_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001011;
  assign _03878_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001010;
  assign _03879_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001001;
  assign _03880_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1001000;
  assign _03881_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000111;
  assign _03882_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000110;
  assign _03883_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000101;
  assign _03884_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000100;
  assign _03885_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000011;
  assign _03886_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000010;
  assign _03887_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000001;
  assign _03888_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 7'b1000000;
  assign _03889_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111111;
  assign _03890_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111110;
  assign _03891_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111101;
  assign _03892_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111100;
  assign _03893_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111011;
  assign _03894_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111010;
  assign _03895_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111001;
  assign _03896_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b111000;
  assign _03897_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110111;
  assign _03898_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110110;
  assign _03899_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110101;
  assign _03900_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110100;
  assign _03901_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110011;
  assign _03902_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110010;
  assign _03903_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110001;
  assign _03904_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b110000;
  assign _03905_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101111;
  assign _03906_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101110;
  assign _03907_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101101;
  assign _03908_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101100;
  assign _03909_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101011;
  assign _03910_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101010;
  assign _03911_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101001;
  assign _03912_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b101000;
  assign _03913_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100111;
  assign _03914_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100110;
  assign _03915_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100101;
  assign _03916_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100100;
  assign _03917_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100011;
  assign _03918_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100010;
  assign _03919_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100001;
  assign _03920_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 6'b100000;
  assign _03921_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11111;
  assign _03922_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11110;
  assign _03923_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11101;
  assign _03924_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11100;
  assign _03925_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11011;
  assign _03926_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11010;
  assign _03927_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11001;
  assign _03928_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b11000;
  assign _03929_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10111;
  assign _03930_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10110;
  assign _03931_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10101;
  assign _03932_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10100;
  assign _03933_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10011;
  assign _03934_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10010;
  assign _03935_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10001;
  assign _03936_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 5'b10000;
  assign _03937_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1111;
  assign _03938_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1110;
  assign _03939_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1101;
  assign _03940_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1100;
  assign _03941_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1011;
  assign _03942_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1010;
  assign _03943_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1001;
  assign _03944_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 4'b1000;
  assign _03945_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 3'b111;
  assign _03946_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 3'b110;
  assign _03947_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 3'b101;
  assign _03948_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 3'b100;
  assign _03949_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 2'b11;
  assign _03950_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 2'b10;
  assign _03951_ = vec_sum_100_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9741" *) 1'b1;
  function [7:0] _13370_;
    input [7:0] a;
    input [799:0] b;
    input [99:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *)
    (* parallel_case *)
    casez (s)
      100'b???????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13370_ = b[7:0];
      100'b??????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13370_ = b[15:8];
      100'b?????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13370_ = b[23:16];
      100'b????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13370_ = b[31:24];
      100'b???????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13370_ = b[39:32];
      100'b??????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13370_ = b[47:40];
      100'b?????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13370_ = b[55:48];
      100'b????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13370_ = b[63:56];
      100'b???????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13370_ = b[71:64];
      100'b??????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13370_ = b[79:72];
      100'b?????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13370_ = b[87:80];
      100'b????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13370_ = b[95:88];
      100'b???????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13370_ = b[103:96];
      100'b??????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13370_ = b[111:104];
      100'b?????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13370_ = b[119:112];
      100'b????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13370_ = b[127:120];
      100'b???????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13370_ = b[135:128];
      100'b??????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13370_ = b[143:136];
      100'b?????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13370_ = b[151:144];
      100'b????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13370_ = b[159:152];
      100'b???????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13370_ = b[167:160];
      100'b??????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13370_ = b[175:168];
      100'b?????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13370_ = b[183:176];
      100'b????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13370_ = b[191:184];
      100'b???????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13370_ = b[199:192];
      100'b??????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13370_ = b[207:200];
      100'b?????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13370_ = b[215:208];
      100'b????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13370_ = b[223:216];
      100'b???????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13370_ = b[231:224];
      100'b??????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13370_ = b[239:232];
      100'b?????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13370_ = b[247:240];
      100'b????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13370_ = b[255:248];
      100'b???????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13370_ = b[263:256];
      100'b??????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13370_ = b[271:264];
      100'b?????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13370_ = b[279:272];
      100'b????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13370_ = b[287:280];
      100'b???????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13370_ = b[295:288];
      100'b??????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13370_ = b[303:296];
      100'b?????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13370_ = b[311:304];
      100'b????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13370_ = b[319:312];
      100'b???????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13370_ = b[327:320];
      100'b??????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13370_ = b[335:328];
      100'b?????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13370_ = b[343:336];
      100'b????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13370_ = b[351:344];
      100'b???????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13370_ = b[359:352];
      100'b??????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13370_ = b[367:360];
      100'b?????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13370_ = b[375:368];
      100'b????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13370_ = b[383:376];
      100'b???????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13370_ = b[391:384];
      100'b??????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13370_ = b[399:392];
      100'b?????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13370_ = b[407:400];
      100'b????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13370_ = b[415:408];
      100'b???????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13370_ = b[423:416];
      100'b??????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13370_ = b[431:424];
      100'b?????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13370_ = b[439:432];
      100'b????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13370_ = b[447:440];
      100'b???????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13370_ = b[455:448];
      100'b??????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13370_ = b[463:456];
      100'b?????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13370_ = b[471:464];
      100'b????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13370_ = b[479:472];
      100'b???????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13370_ = b[487:480];
      100'b??????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13370_ = b[495:488];
      100'b?????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13370_ = b[503:496];
      100'b????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13370_ = b[511:504];
      100'b???????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13370_ = b[519:512];
      100'b??????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13370_ = b[527:520];
      100'b?????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13370_ = b[535:528];
      100'b????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13370_ = b[543:536];
      100'b???????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13370_ = b[551:544];
      100'b??????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13370_ = b[559:552];
      100'b?????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13370_ = b[567:560];
      100'b????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13370_ = b[575:568];
      100'b???????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13370_ = b[583:576];
      100'b??????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13370_ = b[591:584];
      100'b?????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13370_ = b[599:592];
      100'b????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13370_ = b[607:600];
      100'b???????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[615:608];
      100'b??????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[623:616];
      100'b?????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[631:624];
      100'b????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[639:632];
      100'b???????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[647:640];
      100'b??????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[655:648];
      100'b?????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[663:656];
      100'b????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[671:664];
      100'b???????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[679:672];
      100'b??????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[687:680];
      100'b?????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[695:688];
      100'b????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[703:696];
      100'b???????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[711:704];
      100'b??????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[719:712];
      100'b?????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[727:720];
      100'b????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[735:728];
      100'b???????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[743:736];
      100'b??????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[751:744];
      100'b?????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[759:752];
      100'b????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[767:760];
      100'b???1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[775:768];
      100'b??1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[783:776];
      100'b?1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[791:784];
      100'b1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _13370_ = b[799:792];
      default:
        _13370_ = a;
    endcase
  endfunction
  assign vec_data_099 = _13370_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784], data_d1[799:792] }, { _04051_, _04050_, _04049_, _04048_, _04047_, _04046_, _04045_, _04044_, _04043_, _04042_, _04041_, _04040_, _04039_, _04038_, _04037_, _04036_, _04035_, _04034_, _04033_, _04032_, _04031_, _04030_, _04029_, _04028_, _04027_, _04026_, _04025_, _04024_, _04023_, _04022_, _04021_, _04020_, _04019_, _04018_, _04017_, _04016_, _04015_, _04014_, _04013_, _04012_, _04011_, _04010_, _04009_, _04008_, _04007_, _04006_, _04005_, _04004_, _04003_, _04002_, _04001_, _04000_, _03999_, _03998_, _03997_, _03996_, _03995_, _03994_, _03993_, _03992_, _03991_, _03990_, _03989_, _03988_, _03987_, _03986_, _03985_, _03984_, _03983_, _03982_, _03981_, _03980_, _03979_, _03978_, _03977_, _03976_, _03975_, _03974_, _03973_, _03972_, _03971_, _03970_, _03969_, _03968_, _03967_, _03966_, _03965_, _03964_, _03963_, _03962_, _03961_, _03960_, _03959_, _03958_, _03957_, _03956_, _03955_, _03954_, _03953_, _03952_ });
  assign _03952_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1100100;
  assign _03953_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1100011;
  assign _03954_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1100010;
  assign _03955_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1100001;
  assign _03956_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1100000;
  assign _03957_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011111;
  assign _03958_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011110;
  assign _03959_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011101;
  assign _03960_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011100;
  assign _03961_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011011;
  assign _03962_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011010;
  assign _03963_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011001;
  assign _03964_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1011000;
  assign _03965_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010111;
  assign _03966_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010110;
  assign _03967_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010101;
  assign _03968_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010100;
  assign _03969_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010011;
  assign _03970_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010010;
  assign _03971_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010001;
  assign _03972_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1010000;
  assign _03973_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001111;
  assign _03974_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001110;
  assign _03975_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001101;
  assign _03976_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001100;
  assign _03977_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001011;
  assign _03978_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001010;
  assign _03979_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001001;
  assign _03980_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1001000;
  assign _03981_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000111;
  assign _03982_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000110;
  assign _03983_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000101;
  assign _03984_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000100;
  assign _03985_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000011;
  assign _03986_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000010;
  assign _03987_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000001;
  assign _03988_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 7'b1000000;
  assign _03989_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111111;
  assign _03990_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111110;
  assign _03991_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111101;
  assign _03992_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111100;
  assign _03993_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111011;
  assign _03994_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111010;
  assign _03995_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111001;
  assign _03996_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b111000;
  assign _03997_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110111;
  assign _03998_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110110;
  assign _03999_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110101;
  assign _04000_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110100;
  assign _04001_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110011;
  assign _04002_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110010;
  assign _04003_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110001;
  assign _04004_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b110000;
  assign _04005_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101111;
  assign _04006_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101110;
  assign _04007_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101101;
  assign _04008_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101100;
  assign _04009_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101011;
  assign _04010_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101010;
  assign _04011_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101001;
  assign _04012_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b101000;
  assign _04013_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100111;
  assign _04014_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100110;
  assign _04015_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100101;
  assign _04016_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100100;
  assign _04017_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100011;
  assign _04018_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100010;
  assign _04019_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100001;
  assign _04020_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 6'b100000;
  assign _04021_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11111;
  assign _04022_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11110;
  assign _04023_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11101;
  assign _04024_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11100;
  assign _04025_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11011;
  assign _04026_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11010;
  assign _04027_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11001;
  assign _04028_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b11000;
  assign _04029_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10111;
  assign _04030_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10110;
  assign _04031_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10101;
  assign _04032_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10100;
  assign _04033_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10011;
  assign _04034_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10010;
  assign _04035_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10001;
  assign _04036_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 5'b10000;
  assign _04037_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1111;
  assign _04038_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1110;
  assign _04039_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1101;
  assign _04040_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1100;
  assign _04041_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1011;
  assign _04042_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1010;
  assign _04043_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1001;
  assign _04044_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 4'b1000;
  assign _04045_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 3'b111;
  assign _04046_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 3'b110;
  assign _04047_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 3'b101;
  assign _04048_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 3'b100;
  assign _04049_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 2'b11;
  assign _04050_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 2'b10;
  assign _04051_ = vec_sum_099_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9633" *) 1'b1;
  function [7:0] _13471_;
    input [7:0] a;
    input [791:0] b;
    input [98:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *)
    (* parallel_case *)
    casez (s)
      99'b??????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13471_ = b[7:0];
      99'b?????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13471_ = b[15:8];
      99'b????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13471_ = b[23:16];
      99'b???????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13471_ = b[31:24];
      99'b??????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13471_ = b[39:32];
      99'b?????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13471_ = b[47:40];
      99'b????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13471_ = b[55:48];
      99'b???????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13471_ = b[63:56];
      99'b??????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13471_ = b[71:64];
      99'b?????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13471_ = b[79:72];
      99'b????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13471_ = b[87:80];
      99'b???????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13471_ = b[95:88];
      99'b??????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13471_ = b[103:96];
      99'b?????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13471_ = b[111:104];
      99'b????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13471_ = b[119:112];
      99'b???????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13471_ = b[127:120];
      99'b??????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13471_ = b[135:128];
      99'b?????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13471_ = b[143:136];
      99'b????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13471_ = b[151:144];
      99'b???????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13471_ = b[159:152];
      99'b??????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13471_ = b[167:160];
      99'b?????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13471_ = b[175:168];
      99'b????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13471_ = b[183:176];
      99'b???????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13471_ = b[191:184];
      99'b??????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13471_ = b[199:192];
      99'b?????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13471_ = b[207:200];
      99'b????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13471_ = b[215:208];
      99'b???????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13471_ = b[223:216];
      99'b??????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13471_ = b[231:224];
      99'b?????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13471_ = b[239:232];
      99'b????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13471_ = b[247:240];
      99'b???????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13471_ = b[255:248];
      99'b??????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13471_ = b[263:256];
      99'b?????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13471_ = b[271:264];
      99'b????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13471_ = b[279:272];
      99'b???????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13471_ = b[287:280];
      99'b??????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13471_ = b[295:288];
      99'b?????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13471_ = b[303:296];
      99'b????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13471_ = b[311:304];
      99'b???????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13471_ = b[319:312];
      99'b??????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13471_ = b[327:320];
      99'b?????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13471_ = b[335:328];
      99'b????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13471_ = b[343:336];
      99'b???????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13471_ = b[351:344];
      99'b??????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13471_ = b[359:352];
      99'b?????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13471_ = b[367:360];
      99'b????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13471_ = b[375:368];
      99'b???????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13471_ = b[383:376];
      99'b??????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13471_ = b[391:384];
      99'b?????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13471_ = b[399:392];
      99'b????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13471_ = b[407:400];
      99'b???????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13471_ = b[415:408];
      99'b??????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13471_ = b[423:416];
      99'b?????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13471_ = b[431:424];
      99'b????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13471_ = b[439:432];
      99'b???????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13471_ = b[447:440];
      99'b??????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13471_ = b[455:448];
      99'b?????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13471_ = b[463:456];
      99'b????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13471_ = b[471:464];
      99'b???????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13471_ = b[479:472];
      99'b??????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13471_ = b[487:480];
      99'b?????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13471_ = b[495:488];
      99'b????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13471_ = b[503:496];
      99'b???????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13471_ = b[511:504];
      99'b??????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13471_ = b[519:512];
      99'b?????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13471_ = b[527:520];
      99'b????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13471_ = b[535:528];
      99'b???????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13471_ = b[543:536];
      99'b??????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13471_ = b[551:544];
      99'b?????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13471_ = b[559:552];
      99'b????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13471_ = b[567:560];
      99'b???????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13471_ = b[575:568];
      99'b??????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13471_ = b[583:576];
      99'b?????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13471_ = b[591:584];
      99'b????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13471_ = b[599:592];
      99'b???????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13471_ = b[607:600];
      99'b??????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[615:608];
      99'b?????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[623:616];
      99'b????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[631:624];
      99'b???????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[639:632];
      99'b??????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[647:640];
      99'b?????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[655:648];
      99'b????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[663:656];
      99'b???????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[671:664];
      99'b??????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[679:672];
      99'b?????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[687:680];
      99'b????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[695:688];
      99'b???????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[703:696];
      99'b??????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[711:704];
      99'b?????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[719:712];
      99'b????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[727:720];
      99'b???????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[735:728];
      99'b??????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[743:736];
      99'b?????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[751:744];
      99'b????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[759:752];
      99'b???1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[767:760];
      99'b??1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[775:768];
      99'b?1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[783:776];
      99'b1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _13471_ = b[791:784];
      default:
        _13471_ = a;
    endcase
  endfunction
  assign vec_data_098 = _13471_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776], data_d1[791:784] }, { _04150_, _04149_, _04148_, _04147_, _04146_, _04145_, _04144_, _04143_, _04142_, _04141_, _04140_, _04139_, _04138_, _04137_, _04136_, _04135_, _04134_, _04133_, _04132_, _04131_, _04130_, _04129_, _04128_, _04127_, _04126_, _04125_, _04124_, _04123_, _04122_, _04121_, _04120_, _04119_, _04118_, _04117_, _04116_, _04115_, _04114_, _04113_, _04112_, _04111_, _04110_, _04109_, _04108_, _04107_, _04106_, _04105_, _04104_, _04103_, _04102_, _04101_, _04100_, _04099_, _04098_, _04097_, _04096_, _04095_, _04094_, _04093_, _04092_, _04091_, _04090_, _04089_, _04088_, _04087_, _04086_, _04085_, _04084_, _04083_, _04082_, _04081_, _04080_, _04079_, _04078_, _04077_, _04076_, _04075_, _04074_, _04073_, _04072_, _04071_, _04070_, _04069_, _04068_, _04067_, _04066_, _04065_, _04064_, _04063_, _04062_, _04061_, _04060_, _04059_, _04058_, _04057_, _04056_, _04055_, _04054_, _04053_, _04052_ });
  assign _04052_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1100011;
  assign _04053_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1100010;
  assign _04054_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1100001;
  assign _04055_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1100000;
  assign _04056_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011111;
  assign _04057_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011110;
  assign _04058_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011101;
  assign _04059_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011100;
  assign _04060_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011011;
  assign _04061_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011010;
  assign _04062_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011001;
  assign _04063_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1011000;
  assign _04064_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010111;
  assign _04065_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010110;
  assign _04066_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010101;
  assign _04067_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010100;
  assign _04068_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010011;
  assign _04069_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010010;
  assign _04070_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010001;
  assign _04071_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1010000;
  assign _04072_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001111;
  assign _04073_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001110;
  assign _04074_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001101;
  assign _04075_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001100;
  assign _04076_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001011;
  assign _04077_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001010;
  assign _04078_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001001;
  assign _04079_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1001000;
  assign _04080_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000111;
  assign _04081_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000110;
  assign _04082_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000101;
  assign _04083_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000100;
  assign _04084_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000011;
  assign _04085_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000010;
  assign _04086_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000001;
  assign _04087_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 7'b1000000;
  assign _04088_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111111;
  assign _04089_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111110;
  assign _04090_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111101;
  assign _04091_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111100;
  assign _04092_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111011;
  assign _04093_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111010;
  assign _04094_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111001;
  assign _04095_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b111000;
  assign _04096_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110111;
  assign _04097_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110110;
  assign _04098_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110101;
  assign _04099_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110100;
  assign _04100_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110011;
  assign _04101_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110010;
  assign _04102_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110001;
  assign _04103_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b110000;
  assign _04104_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101111;
  assign _04105_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101110;
  assign _04106_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101101;
  assign _04107_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101100;
  assign _04108_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101011;
  assign _04109_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101010;
  assign _04110_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101001;
  assign _04111_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b101000;
  assign _04112_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100111;
  assign _04113_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100110;
  assign _04114_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100101;
  assign _04115_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100100;
  assign _04116_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100011;
  assign _04117_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100010;
  assign _04118_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100001;
  assign _04119_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 6'b100000;
  assign _04120_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11111;
  assign _04121_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11110;
  assign _04122_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11101;
  assign _04123_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11100;
  assign _04124_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11011;
  assign _04125_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11010;
  assign _04126_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11001;
  assign _04127_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b11000;
  assign _04128_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10111;
  assign _04129_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10110;
  assign _04130_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10101;
  assign _04131_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10100;
  assign _04132_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10011;
  assign _04133_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10010;
  assign _04134_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10001;
  assign _04135_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 5'b10000;
  assign _04136_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1111;
  assign _04137_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1110;
  assign _04138_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1101;
  assign _04139_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1100;
  assign _04140_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1011;
  assign _04141_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1010;
  assign _04142_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1001;
  assign _04143_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 4'b1000;
  assign _04144_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 3'b111;
  assign _04145_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 3'b110;
  assign _04146_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 3'b101;
  assign _04147_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 3'b100;
  assign _04148_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 2'b11;
  assign _04149_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 2'b10;
  assign _04150_ = vec_sum_098_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9526" *) 1'b1;
  function [7:0] _13571_;
    input [7:0] a;
    input [783:0] b;
    input [97:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *)
    (* parallel_case *)
    casez (s)
      98'b?????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13571_ = b[7:0];
      98'b????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13571_ = b[15:8];
      98'b???????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13571_ = b[23:16];
      98'b??????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13571_ = b[31:24];
      98'b?????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13571_ = b[39:32];
      98'b????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13571_ = b[47:40];
      98'b???????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13571_ = b[55:48];
      98'b??????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13571_ = b[63:56];
      98'b?????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13571_ = b[71:64];
      98'b????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13571_ = b[79:72];
      98'b???????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13571_ = b[87:80];
      98'b??????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13571_ = b[95:88];
      98'b?????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13571_ = b[103:96];
      98'b????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13571_ = b[111:104];
      98'b???????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13571_ = b[119:112];
      98'b??????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13571_ = b[127:120];
      98'b?????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13571_ = b[135:128];
      98'b????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13571_ = b[143:136];
      98'b???????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13571_ = b[151:144];
      98'b??????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13571_ = b[159:152];
      98'b?????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13571_ = b[167:160];
      98'b????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13571_ = b[175:168];
      98'b???????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13571_ = b[183:176];
      98'b??????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13571_ = b[191:184];
      98'b?????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13571_ = b[199:192];
      98'b????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13571_ = b[207:200];
      98'b???????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13571_ = b[215:208];
      98'b??????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13571_ = b[223:216];
      98'b?????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13571_ = b[231:224];
      98'b????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13571_ = b[239:232];
      98'b???????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13571_ = b[247:240];
      98'b??????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13571_ = b[255:248];
      98'b?????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13571_ = b[263:256];
      98'b????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13571_ = b[271:264];
      98'b???????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13571_ = b[279:272];
      98'b??????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13571_ = b[287:280];
      98'b?????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13571_ = b[295:288];
      98'b????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13571_ = b[303:296];
      98'b???????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13571_ = b[311:304];
      98'b??????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13571_ = b[319:312];
      98'b?????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13571_ = b[327:320];
      98'b????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13571_ = b[335:328];
      98'b???????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13571_ = b[343:336];
      98'b??????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13571_ = b[351:344];
      98'b?????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13571_ = b[359:352];
      98'b????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13571_ = b[367:360];
      98'b???????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13571_ = b[375:368];
      98'b??????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13571_ = b[383:376];
      98'b?????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13571_ = b[391:384];
      98'b????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13571_ = b[399:392];
      98'b???????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13571_ = b[407:400];
      98'b??????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13571_ = b[415:408];
      98'b?????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13571_ = b[423:416];
      98'b????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13571_ = b[431:424];
      98'b???????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13571_ = b[439:432];
      98'b??????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13571_ = b[447:440];
      98'b?????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13571_ = b[455:448];
      98'b????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13571_ = b[463:456];
      98'b???????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13571_ = b[471:464];
      98'b??????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13571_ = b[479:472];
      98'b?????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13571_ = b[487:480];
      98'b????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13571_ = b[495:488];
      98'b???????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13571_ = b[503:496];
      98'b??????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13571_ = b[511:504];
      98'b?????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13571_ = b[519:512];
      98'b????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13571_ = b[527:520];
      98'b???????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13571_ = b[535:528];
      98'b??????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13571_ = b[543:536];
      98'b?????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13571_ = b[551:544];
      98'b????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13571_ = b[559:552];
      98'b???????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13571_ = b[567:560];
      98'b??????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13571_ = b[575:568];
      98'b?????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13571_ = b[583:576];
      98'b????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13571_ = b[591:584];
      98'b???????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13571_ = b[599:592];
      98'b??????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13571_ = b[607:600];
      98'b?????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[615:608];
      98'b????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[623:616];
      98'b???????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[631:624];
      98'b??????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[639:632];
      98'b?????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[647:640];
      98'b????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[655:648];
      98'b???????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[663:656];
      98'b??????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[671:664];
      98'b?????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[679:672];
      98'b????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[687:680];
      98'b???????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[695:688];
      98'b??????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[703:696];
      98'b?????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[711:704];
      98'b????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[719:712];
      98'b???????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[727:720];
      98'b??????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[735:728];
      98'b?????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[743:736];
      98'b????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[751:744];
      98'b???1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[759:752];
      98'b??1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[767:760];
      98'b?1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[775:768];
      98'b1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _13571_ = b[783:776];
      default:
        _13571_ = a;
    endcase
  endfunction
  assign vec_data_097 = _13571_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768], data_d1[783:776] }, { _04248_, _04247_, _04246_, _04245_, _04244_, _04243_, _04242_, _04241_, _04240_, _04239_, _04238_, _04237_, _04236_, _04235_, _04234_, _04233_, _04232_, _04231_, _04230_, _04229_, _04228_, _04227_, _04226_, _04225_, _04224_, _04223_, _04222_, _04221_, _04220_, _04219_, _04218_, _04217_, _04216_, _04215_, _04214_, _04213_, _04212_, _04211_, _04210_, _04209_, _04208_, _04207_, _04206_, _04205_, _04204_, _04203_, _04202_, _04201_, _04200_, _04199_, _04198_, _04197_, _04196_, _04195_, _04194_, _04193_, _04192_, _04191_, _04190_, _04189_, _04188_, _04187_, _04186_, _04185_, _04184_, _04183_, _04182_, _04181_, _04180_, _04179_, _04178_, _04177_, _04176_, _04175_, _04174_, _04173_, _04172_, _04171_, _04170_, _04169_, _04168_, _04167_, _04166_, _04165_, _04164_, _04163_, _04162_, _04161_, _04160_, _04159_, _04158_, _04157_, _04156_, _04155_, _04154_, _04153_, _04152_, _04151_ });
  assign _04151_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1100010;
  assign _04152_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1100001;
  assign _04153_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1100000;
  assign _04154_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011111;
  assign _04155_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011110;
  assign _04156_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011101;
  assign _04157_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011100;
  assign _04158_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011011;
  assign _04159_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011010;
  assign _04160_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011001;
  assign _04161_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1011000;
  assign _04162_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010111;
  assign _04163_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010110;
  assign _04164_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010101;
  assign _04165_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010100;
  assign _04166_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010011;
  assign _04167_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010010;
  assign _04168_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010001;
  assign _04169_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1010000;
  assign _04170_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001111;
  assign _04171_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001110;
  assign _04172_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001101;
  assign _04173_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001100;
  assign _04174_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001011;
  assign _04175_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001010;
  assign _04176_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001001;
  assign _04177_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1001000;
  assign _04178_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000111;
  assign _04179_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000110;
  assign _04180_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000101;
  assign _04181_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000100;
  assign _04182_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000011;
  assign _04183_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000010;
  assign _04184_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000001;
  assign _04185_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 7'b1000000;
  assign _04186_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111111;
  assign _04187_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111110;
  assign _04188_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111101;
  assign _04189_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111100;
  assign _04190_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111011;
  assign _04191_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111010;
  assign _04192_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111001;
  assign _04193_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b111000;
  assign _04194_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110111;
  assign _04195_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110110;
  assign _04196_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110101;
  assign _04197_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110100;
  assign _04198_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110011;
  assign _04199_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110010;
  assign _04200_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110001;
  assign _04201_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b110000;
  assign _04202_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101111;
  assign _04203_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101110;
  assign _04204_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101101;
  assign _04205_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101100;
  assign _04206_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101011;
  assign _04207_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101010;
  assign _04208_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101001;
  assign _04209_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b101000;
  assign _04210_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100111;
  assign _04211_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100110;
  assign _04212_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100101;
  assign _04213_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100100;
  assign _04214_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100011;
  assign _04215_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100010;
  assign _04216_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100001;
  assign _04217_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 6'b100000;
  assign _04218_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11111;
  assign _04219_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11110;
  assign _04220_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11101;
  assign _04221_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11100;
  assign _04222_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11011;
  assign _04223_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11010;
  assign _04224_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11001;
  assign _04225_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b11000;
  assign _04226_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10111;
  assign _04227_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10110;
  assign _04228_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10101;
  assign _04229_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10100;
  assign _04230_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10011;
  assign _04231_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10010;
  assign _04232_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10001;
  assign _04233_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 5'b10000;
  assign _04234_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1111;
  assign _04235_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1110;
  assign _04236_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1101;
  assign _04237_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1100;
  assign _04238_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1011;
  assign _04239_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1010;
  assign _04240_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1001;
  assign _04241_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 4'b1000;
  assign _04242_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 3'b111;
  assign _04243_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 3'b110;
  assign _04244_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 3'b101;
  assign _04245_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 3'b100;
  assign _04246_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 2'b11;
  assign _04247_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 2'b10;
  assign _04248_ = vec_sum_097_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9420" *) 1'b1;
  function [7:0] _13670_;
    input [7:0] a;
    input [775:0] b;
    input [96:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *)
    (* parallel_case *)
    casez (s)
      97'b????????????????????????????????????????????????????????????????????????????????????????????????1:
        _13670_ = b[7:0];
      97'b???????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13670_ = b[15:8];
      97'b??????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13670_ = b[23:16];
      97'b?????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13670_ = b[31:24];
      97'b????????????????????????????????????????????????????????????????????????????????????????????1????:
        _13670_ = b[39:32];
      97'b???????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13670_ = b[47:40];
      97'b??????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13670_ = b[55:48];
      97'b?????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13670_ = b[63:56];
      97'b????????????????????????????????????????????????????????????????????????????????????????1????????:
        _13670_ = b[71:64];
      97'b???????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13670_ = b[79:72];
      97'b??????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13670_ = b[87:80];
      97'b?????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13670_ = b[95:88];
      97'b????????????????????????????????????????????????????????????????????????????????????1????????????:
        _13670_ = b[103:96];
      97'b???????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13670_ = b[111:104];
      97'b??????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13670_ = b[119:112];
      97'b?????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13670_ = b[127:120];
      97'b????????????????????????????????????????????????????????????????????????????????1????????????????:
        _13670_ = b[135:128];
      97'b???????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13670_ = b[143:136];
      97'b??????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13670_ = b[151:144];
      97'b?????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13670_ = b[159:152];
      97'b????????????????????????????????????????????????????????????????????????????1????????????????????:
        _13670_ = b[167:160];
      97'b???????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13670_ = b[175:168];
      97'b??????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13670_ = b[183:176];
      97'b?????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13670_ = b[191:184];
      97'b????????????????????????????????????????????????????????????????????????1????????????????????????:
        _13670_ = b[199:192];
      97'b???????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13670_ = b[207:200];
      97'b??????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13670_ = b[215:208];
      97'b?????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13670_ = b[223:216];
      97'b????????????????????????????????????????????????????????????????????1????????????????????????????:
        _13670_ = b[231:224];
      97'b???????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13670_ = b[239:232];
      97'b??????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13670_ = b[247:240];
      97'b?????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13670_ = b[255:248];
      97'b????????????????????????????????????????????????????????????????1????????????????????????????????:
        _13670_ = b[263:256];
      97'b???????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13670_ = b[271:264];
      97'b??????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13670_ = b[279:272];
      97'b?????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13670_ = b[287:280];
      97'b????????????????????????????????????????????????????????????1????????????????????????????????????:
        _13670_ = b[295:288];
      97'b???????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13670_ = b[303:296];
      97'b??????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13670_ = b[311:304];
      97'b?????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13670_ = b[319:312];
      97'b????????????????????????????????????????????????????????1????????????????????????????????????????:
        _13670_ = b[327:320];
      97'b???????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13670_ = b[335:328];
      97'b??????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13670_ = b[343:336];
      97'b?????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13670_ = b[351:344];
      97'b????????????????????????????????????????????????????1????????????????????????????????????????????:
        _13670_ = b[359:352];
      97'b???????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13670_ = b[367:360];
      97'b??????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13670_ = b[375:368];
      97'b?????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13670_ = b[383:376];
      97'b????????????????????????????????????????????????1????????????????????????????????????????????????:
        _13670_ = b[391:384];
      97'b???????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13670_ = b[399:392];
      97'b??????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13670_ = b[407:400];
      97'b?????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13670_ = b[415:408];
      97'b????????????????????????????????????????????1????????????????????????????????????????????????????:
        _13670_ = b[423:416];
      97'b???????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13670_ = b[431:424];
      97'b??????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13670_ = b[439:432];
      97'b?????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13670_ = b[447:440];
      97'b????????????????????????????????????????1????????????????????????????????????????????????????????:
        _13670_ = b[455:448];
      97'b???????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13670_ = b[463:456];
      97'b??????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13670_ = b[471:464];
      97'b?????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13670_ = b[479:472];
      97'b????????????????????????????????????1????????????????????????????????????????????????????????????:
        _13670_ = b[487:480];
      97'b???????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13670_ = b[495:488];
      97'b??????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13670_ = b[503:496];
      97'b?????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13670_ = b[511:504];
      97'b????????????????????????????????1????????????????????????????????????????????????????????????????:
        _13670_ = b[519:512];
      97'b???????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13670_ = b[527:520];
      97'b??????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13670_ = b[535:528];
      97'b?????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13670_ = b[543:536];
      97'b????????????????????????????1????????????????????????????????????????????????????????????????????:
        _13670_ = b[551:544];
      97'b???????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13670_ = b[559:552];
      97'b??????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13670_ = b[567:560];
      97'b?????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13670_ = b[575:568];
      97'b????????????????????????1????????????????????????????????????????????????????????????????????????:
        _13670_ = b[583:576];
      97'b???????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13670_ = b[591:584];
      97'b??????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13670_ = b[599:592];
      97'b?????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13670_ = b[607:600];
      97'b????????????????????1????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[615:608];
      97'b???????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[623:616];
      97'b??????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[631:624];
      97'b?????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[639:632];
      97'b????????????????1????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[647:640];
      97'b???????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[655:648];
      97'b??????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[663:656];
      97'b?????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[671:664];
      97'b????????????1????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[679:672];
      97'b???????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[687:680];
      97'b??????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[695:688];
      97'b?????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[703:696];
      97'b????????1????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[711:704];
      97'b???????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[719:712];
      97'b??????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[727:720];
      97'b?????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[735:728];
      97'b????1????????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[743:736];
      97'b???1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[751:744];
      97'b??1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[759:752];
      97'b?1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[767:760];
      97'b1????????????????????????????????????????????????????????????????????????????????????????????????:
        _13670_ = b[775:768];
      default:
        _13670_ = a;
    endcase
  endfunction
  assign vec_data_096 = _13670_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760], data_d1[775:768] }, { _04345_, _04344_, _04343_, _04342_, _04341_, _04340_, _04339_, _04338_, _04337_, _04336_, _04335_, _04334_, _04333_, _04332_, _04331_, _04330_, _04329_, _04328_, _04327_, _04326_, _04325_, _04324_, _04323_, _04322_, _04321_, _04320_, _04319_, _04318_, _04317_, _04316_, _04315_, _04314_, _04313_, _04312_, _04311_, _04310_, _04309_, _04308_, _04307_, _04306_, _04305_, _04304_, _04303_, _04302_, _04301_, _04300_, _04299_, _04298_, _04297_, _04296_, _04295_, _04294_, _04293_, _04292_, _04291_, _04290_, _04289_, _04288_, _04287_, _04286_, _04285_, _04284_, _04283_, _04282_, _04281_, _04280_, _04279_, _04278_, _04277_, _04276_, _04275_, _04274_, _04273_, _04272_, _04271_, _04270_, _04269_, _04268_, _04267_, _04266_, _04265_, _04264_, _04263_, _04262_, _04261_, _04260_, _04259_, _04258_, _04257_, _04256_, _04255_, _04254_, _04253_, _04252_, _04251_, _04250_, _04249_ });
  assign _04249_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1100001;
  assign _04250_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1100000;
  assign _04251_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9410|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011111;
  assign _04252_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9409|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011110;
  assign _04253_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011101;
  assign _04254_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011100;
  assign _04255_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011011;
  assign _04256_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011010;
  assign _04257_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011001;
  assign _04258_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1011000;
  assign _04259_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010111;
  assign _04260_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010110;
  assign _04261_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010101;
  assign _04262_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010100;
  assign _04263_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010011;
  assign _04264_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010010;
  assign _04265_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010001;
  assign _04266_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1010000;
  assign _04267_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001111;
  assign _04268_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001110;
  assign _04269_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001101;
  assign _04270_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001100;
  assign _04271_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001011;
  assign _04272_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001010;
  assign _04273_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001001;
  assign _04274_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1001000;
  assign _04275_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000111;
  assign _04276_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000110;
  assign _04277_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000101;
  assign _04278_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000100;
  assign _04279_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000011;
  assign _04280_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000010;
  assign _04281_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000001;
  assign _04282_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 7'b1000000;
  assign _04283_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111111;
  assign _04284_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111110;
  assign _04285_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111101;
  assign _04286_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111100;
  assign _04287_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111011;
  assign _04288_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111010;
  assign _04289_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111001;
  assign _04290_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b111000;
  assign _04291_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110111;
  assign _04292_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110110;
  assign _04293_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110101;
  assign _04294_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110100;
  assign _04295_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110011;
  assign _04296_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110010;
  assign _04297_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110001;
  assign _04298_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b110000;
  assign _04299_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101111;
  assign _04300_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101110;
  assign _04301_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101101;
  assign _04302_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101100;
  assign _04303_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101011;
  assign _04304_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101010;
  assign _04305_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101001;
  assign _04306_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b101000;
  assign _04307_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100111;
  assign _04308_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100110;
  assign _04309_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100101;
  assign _04310_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100100;
  assign _04311_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100011;
  assign _04312_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100010;
  assign _04313_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100001;
  assign _04314_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 6'b100000;
  assign _04315_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11111;
  assign _04316_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11110;
  assign _04317_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11101;
  assign _04318_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11100;
  assign _04319_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11011;
  assign _04320_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11010;
  assign _04321_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11001;
  assign _04322_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b11000;
  assign _04323_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10111;
  assign _04324_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10110;
  assign _04325_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10101;
  assign _04326_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10100;
  assign _04327_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10011;
  assign _04328_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10010;
  assign _04329_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10001;
  assign _04330_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 5'b10000;
  assign _04331_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1111;
  assign _04332_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1110;
  assign _04333_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1101;
  assign _04334_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1100;
  assign _04335_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1011;
  assign _04336_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1010;
  assign _04337_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1001;
  assign _04338_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 4'b1000;
  assign _04339_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 3'b111;
  assign _04340_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 3'b110;
  assign _04341_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 3'b101;
  assign _04342_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 3'b100;
  assign _04343_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 2'b11;
  assign _04344_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 2'b10;
  assign _04345_ = vec_sum_096_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9315" *) 1'b1;
  function [7:0] _13768_;
    input [7:0] a;
    input [767:0] b;
    input [95:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *)
    (* parallel_case *)
    casez (s)
      96'b???????????????????????????????????????????????????????????????????????????????????????????????1:
        _13768_ = b[7:0];
      96'b??????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13768_ = b[15:8];
      96'b?????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13768_ = b[23:16];
      96'b????????????????????????????????????????????????????????????????????????????????????????????1???:
        _13768_ = b[31:24];
      96'b???????????????????????????????????????????????????????????????????????????????????????????1????:
        _13768_ = b[39:32];
      96'b??????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13768_ = b[47:40];
      96'b?????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13768_ = b[55:48];
      96'b????????????????????????????????????????????????????????????????????????????????????????1???????:
        _13768_ = b[63:56];
      96'b???????????????????????????????????????????????????????????????????????????????????????1????????:
        _13768_ = b[71:64];
      96'b??????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13768_ = b[79:72];
      96'b?????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13768_ = b[87:80];
      96'b????????????????????????????????????????????????????????????????????????????????????1???????????:
        _13768_ = b[95:88];
      96'b???????????????????????????????????????????????????????????????????????????????????1????????????:
        _13768_ = b[103:96];
      96'b??????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13768_ = b[111:104];
      96'b?????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13768_ = b[119:112];
      96'b????????????????????????????????????????????????????????????????????????????????1???????????????:
        _13768_ = b[127:120];
      96'b???????????????????????????????????????????????????????????????????????????????1????????????????:
        _13768_ = b[135:128];
      96'b??????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13768_ = b[143:136];
      96'b?????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13768_ = b[151:144];
      96'b????????????????????????????????????????????????????????????????????????????1???????????????????:
        _13768_ = b[159:152];
      96'b???????????????????????????????????????????????????????????????????????????1????????????????????:
        _13768_ = b[167:160];
      96'b??????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13768_ = b[175:168];
      96'b?????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13768_ = b[183:176];
      96'b????????????????????????????????????????????????????????????????????????1???????????????????????:
        _13768_ = b[191:184];
      96'b???????????????????????????????????????????????????????????????????????1????????????????????????:
        _13768_ = b[199:192];
      96'b??????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13768_ = b[207:200];
      96'b?????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13768_ = b[215:208];
      96'b????????????????????????????????????????????????????????????????????1???????????????????????????:
        _13768_ = b[223:216];
      96'b???????????????????????????????????????????????????????????????????1????????????????????????????:
        _13768_ = b[231:224];
      96'b??????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13768_ = b[239:232];
      96'b?????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13768_ = b[247:240];
      96'b????????????????????????????????????????????????????????????????1???????????????????????????????:
        _13768_ = b[255:248];
      96'b???????????????????????????????????????????????????????????????1????????????????????????????????:
        _13768_ = b[263:256];
      96'b??????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13768_ = b[271:264];
      96'b?????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13768_ = b[279:272];
      96'b????????????????????????????????????????????????????????????1???????????????????????????????????:
        _13768_ = b[287:280];
      96'b???????????????????????????????????????????????????????????1????????????????????????????????????:
        _13768_ = b[295:288];
      96'b??????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13768_ = b[303:296];
      96'b?????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13768_ = b[311:304];
      96'b????????????????????????????????????????????????????????1???????????????????????????????????????:
        _13768_ = b[319:312];
      96'b???????????????????????????????????????????????????????1????????????????????????????????????????:
        _13768_ = b[327:320];
      96'b??????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13768_ = b[335:328];
      96'b?????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13768_ = b[343:336];
      96'b????????????????????????????????????????????????????1???????????????????????????????????????????:
        _13768_ = b[351:344];
      96'b???????????????????????????????????????????????????1????????????????????????????????????????????:
        _13768_ = b[359:352];
      96'b??????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13768_ = b[367:360];
      96'b?????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13768_ = b[375:368];
      96'b????????????????????????????????????????????????1???????????????????????????????????????????????:
        _13768_ = b[383:376];
      96'b???????????????????????????????????????????????1????????????????????????????????????????????????:
        _13768_ = b[391:384];
      96'b??????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13768_ = b[399:392];
      96'b?????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13768_ = b[407:400];
      96'b????????????????????????????????????????????1???????????????????????????????????????????????????:
        _13768_ = b[415:408];
      96'b???????????????????????????????????????????1????????????????????????????????????????????????????:
        _13768_ = b[423:416];
      96'b??????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13768_ = b[431:424];
      96'b?????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13768_ = b[439:432];
      96'b????????????????????????????????????????1???????????????????????????????????????????????????????:
        _13768_ = b[447:440];
      96'b???????????????????????????????????????1????????????????????????????????????????????????????????:
        _13768_ = b[455:448];
      96'b??????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13768_ = b[463:456];
      96'b?????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13768_ = b[471:464];
      96'b????????????????????????????????????1???????????????????????????????????????????????????????????:
        _13768_ = b[479:472];
      96'b???????????????????????????????????1????????????????????????????????????????????????????????????:
        _13768_ = b[487:480];
      96'b??????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13768_ = b[495:488];
      96'b?????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13768_ = b[503:496];
      96'b????????????????????????????????1???????????????????????????????????????????????????????????????:
        _13768_ = b[511:504];
      96'b???????????????????????????????1????????????????????????????????????????????????????????????????:
        _13768_ = b[519:512];
      96'b??????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13768_ = b[527:520];
      96'b?????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13768_ = b[535:528];
      96'b????????????????????????????1???????????????????????????????????????????????????????????????????:
        _13768_ = b[543:536];
      96'b???????????????????????????1????????????????????????????????????????????????????????????????????:
        _13768_ = b[551:544];
      96'b??????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13768_ = b[559:552];
      96'b?????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13768_ = b[567:560];
      96'b????????????????????????1???????????????????????????????????????????????????????????????????????:
        _13768_ = b[575:568];
      96'b???????????????????????1????????????????????????????????????????????????????????????????????????:
        _13768_ = b[583:576];
      96'b??????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13768_ = b[591:584];
      96'b?????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13768_ = b[599:592];
      96'b????????????????????1???????????????????????????????????????????????????????????????????????????:
        _13768_ = b[607:600];
      96'b???????????????????1????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[615:608];
      96'b??????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[623:616];
      96'b?????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[631:624];
      96'b????????????????1???????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[639:632];
      96'b???????????????1????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[647:640];
      96'b??????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[655:648];
      96'b?????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[663:656];
      96'b????????????1???????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[671:664];
      96'b???????????1????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[679:672];
      96'b??????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[687:680];
      96'b?????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[695:688];
      96'b????????1???????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[703:696];
      96'b???????1????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[711:704];
      96'b??????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[719:712];
      96'b?????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[727:720];
      96'b????1???????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[735:728];
      96'b???1????????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[743:736];
      96'b??1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[751:744];
      96'b?1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[759:752];
      96'b1???????????????????????????????????????????????????????????????????????????????????????????????:
        _13768_ = b[767:760];
      default:
        _13768_ = a;
    endcase
  endfunction
  assign vec_data_095 = _13768_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752], data_d1[767:760] }, { _04441_, _04440_, _04439_, _04438_, _04437_, _04436_, _04435_, _04434_, _04433_, _04432_, _04431_, _04430_, _04429_, _04428_, _04427_, _04426_, _04425_, _04424_, _04423_, _04422_, _04421_, _04420_, _04419_, _04418_, _04417_, _04416_, _04415_, _04414_, _04413_, _04412_, _04411_, _04410_, _04409_, _04408_, _04407_, _04406_, _04405_, _04404_, _04403_, _04402_, _04401_, _04400_, _04399_, _04398_, _04397_, _04396_, _04395_, _04394_, _04393_, _04392_, _04391_, _04390_, _04389_, _04388_, _04387_, _04386_, _04385_, _04384_, _04383_, _04382_, _04381_, _04380_, _04379_, _04378_, _04377_, _04376_, _04375_, _04374_, _04373_, _04372_, _04371_, _04370_, _04369_, _04368_, _04367_, _04366_, _04365_, _04364_, _04363_, _04362_, _04361_, _04360_, _04359_, _04358_, _04357_, _04356_, _04355_, _04354_, _04353_, _04352_, _04351_, _04350_, _04349_, _04348_, _04347_, _04346_ });
  assign _04346_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1100000;
  assign _04347_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011111;
  assign _04348_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011110;
  assign _04349_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011101;
  assign _04350_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011100;
  assign _04351_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011011;
  assign _04352_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011010;
  assign _04353_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011001;
  assign _04354_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1011000;
  assign _04355_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010111;
  assign _04356_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010110;
  assign _04357_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010101;
  assign _04358_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010100;
  assign _04359_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010011;
  assign _04360_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010010;
  assign _04361_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010001;
  assign _04362_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1010000;
  assign _04363_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001111;
  assign _04364_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001110;
  assign _04365_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001101;
  assign _04366_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001100;
  assign _04367_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001011;
  assign _04368_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001010;
  assign _04369_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001001;
  assign _04370_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1001000;
  assign _04371_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000111;
  assign _04372_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000110;
  assign _04373_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000101;
  assign _04374_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000100;
  assign _04375_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000011;
  assign _04376_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000010;
  assign _04377_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000001;
  assign _04378_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 7'b1000000;
  assign _04379_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111111;
  assign _04380_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111110;
  assign _04381_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111101;
  assign _04382_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111100;
  assign _04383_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111011;
  assign _04384_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111010;
  assign _04385_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111001;
  assign _04386_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b111000;
  assign _04387_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110111;
  assign _04388_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110110;
  assign _04389_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110101;
  assign _04390_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110100;
  assign _04391_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110011;
  assign _04392_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110010;
  assign _04393_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110001;
  assign _04394_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b110000;
  assign _04395_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101111;
  assign _04396_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101110;
  assign _04397_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101101;
  assign _04398_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101100;
  assign _04399_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101011;
  assign _04400_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101010;
  assign _04401_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101001;
  assign _04402_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b101000;
  assign _04403_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100111;
  assign _04404_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100110;
  assign _04405_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100101;
  assign _04406_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100100;
  assign _04407_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100011;
  assign _04408_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100010;
  assign _04409_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100001;
  assign _04410_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 6'b100000;
  assign _04411_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11111;
  assign _04412_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11110;
  assign _04413_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11101;
  assign _04414_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11100;
  assign _04415_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11011;
  assign _04416_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11010;
  assign _04417_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11001;
  assign _04418_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b11000;
  assign _04419_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10111;
  assign _04420_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9233|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10110;
  assign _04421_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10101;
  assign _04422_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10100;
  assign _04423_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10011;
  assign _04424_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10010;
  assign _04425_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10001;
  assign _04426_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 5'b10000;
  assign _04427_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1111;
  assign _04428_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1110;
  assign _04429_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1101;
  assign _04430_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1100;
  assign _04431_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1011;
  assign _04432_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1010;
  assign _04433_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1001;
  assign _04434_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 4'b1000;
  assign _04435_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 3'b111;
  assign _04436_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 3'b110;
  assign _04437_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 3'b101;
  assign _04438_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 3'b100;
  assign _04439_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 2'b11;
  assign _04440_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 2'b10;
  assign _04441_ = vec_sum_095_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9211" *) 1'b1;
  function [7:0] _13865_;
    input [7:0] a;
    input [759:0] b;
    input [94:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *)
    (* parallel_case *)
    casez (s)
      95'b??????????????????????????????????????????????????????????????????????????????????????????????1:
        _13865_ = b[7:0];
      95'b?????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13865_ = b[15:8];
      95'b????????????????????????????????????????????????????????????????????????????????????????????1??:
        _13865_ = b[23:16];
      95'b???????????????????????????????????????????????????????????????????????????????????????????1???:
        _13865_ = b[31:24];
      95'b??????????????????????????????????????????????????????????????????????????????????????????1????:
        _13865_ = b[39:32];
      95'b?????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13865_ = b[47:40];
      95'b????????????????????????????????????????????????????????????????????????????????????????1??????:
        _13865_ = b[55:48];
      95'b???????????????????????????????????????????????????????????????????????????????????????1???????:
        _13865_ = b[63:56];
      95'b??????????????????????????????????????????????????????????????????????????????????????1????????:
        _13865_ = b[71:64];
      95'b?????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13865_ = b[79:72];
      95'b????????????????????????????????????????????????????????????????????????????????????1??????????:
        _13865_ = b[87:80];
      95'b???????????????????????????????????????????????????????????????????????????????????1???????????:
        _13865_ = b[95:88];
      95'b??????????????????????????????????????????????????????????????????????????????????1????????????:
        _13865_ = b[103:96];
      95'b?????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13865_ = b[111:104];
      95'b????????????????????????????????????????????????????????????????????????????????1??????????????:
        _13865_ = b[119:112];
      95'b???????????????????????????????????????????????????????????????????????????????1???????????????:
        _13865_ = b[127:120];
      95'b??????????????????????????????????????????????????????????????????????????????1????????????????:
        _13865_ = b[135:128];
      95'b?????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13865_ = b[143:136];
      95'b????????????????????????????????????????????????????????????????????????????1??????????????????:
        _13865_ = b[151:144];
      95'b???????????????????????????????????????????????????????????????????????????1???????????????????:
        _13865_ = b[159:152];
      95'b??????????????????????????????????????????????????????????????????????????1????????????????????:
        _13865_ = b[167:160];
      95'b?????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13865_ = b[175:168];
      95'b????????????????????????????????????????????????????????????????????????1??????????????????????:
        _13865_ = b[183:176];
      95'b???????????????????????????????????????????????????????????????????????1???????????????????????:
        _13865_ = b[191:184];
      95'b??????????????????????????????????????????????????????????????????????1????????????????????????:
        _13865_ = b[199:192];
      95'b?????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13865_ = b[207:200];
      95'b????????????????????????????????????????????????????????????????????1??????????????????????????:
        _13865_ = b[215:208];
      95'b???????????????????????????????????????????????????????????????????1???????????????????????????:
        _13865_ = b[223:216];
      95'b??????????????????????????????????????????????????????????????????1????????????????????????????:
        _13865_ = b[231:224];
      95'b?????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13865_ = b[239:232];
      95'b????????????????????????????????????????????????????????????????1??????????????????????????????:
        _13865_ = b[247:240];
      95'b???????????????????????????????????????????????????????????????1???????????????????????????????:
        _13865_ = b[255:248];
      95'b??????????????????????????????????????????????????????????????1????????????????????????????????:
        _13865_ = b[263:256];
      95'b?????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13865_ = b[271:264];
      95'b????????????????????????????????????????????????????????????1??????????????????????????????????:
        _13865_ = b[279:272];
      95'b???????????????????????????????????????????????????????????1???????????????????????????????????:
        _13865_ = b[287:280];
      95'b??????????????????????????????????????????????????????????1????????????????????????????????????:
        _13865_ = b[295:288];
      95'b?????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13865_ = b[303:296];
      95'b????????????????????????????????????????????????????????1??????????????????????????????????????:
        _13865_ = b[311:304];
      95'b???????????????????????????????????????????????????????1???????????????????????????????????????:
        _13865_ = b[319:312];
      95'b??????????????????????????????????????????????????????1????????????????????????????????????????:
        _13865_ = b[327:320];
      95'b?????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13865_ = b[335:328];
      95'b????????????????????????????????????????????????????1??????????????????????????????????????????:
        _13865_ = b[343:336];
      95'b???????????????????????????????????????????????????1???????????????????????????????????????????:
        _13865_ = b[351:344];
      95'b??????????????????????????????????????????????????1????????????????????????????????????????????:
        _13865_ = b[359:352];
      95'b?????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13865_ = b[367:360];
      95'b????????????????????????????????????????????????1??????????????????????????????????????????????:
        _13865_ = b[375:368];
      95'b???????????????????????????????????????????????1???????????????????????????????????????????????:
        _13865_ = b[383:376];
      95'b??????????????????????????????????????????????1????????????????????????????????????????????????:
        _13865_ = b[391:384];
      95'b?????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13865_ = b[399:392];
      95'b????????????????????????????????????????????1??????????????????????????????????????????????????:
        _13865_ = b[407:400];
      95'b???????????????????????????????????????????1???????????????????????????????????????????????????:
        _13865_ = b[415:408];
      95'b??????????????????????????????????????????1????????????????????????????????????????????????????:
        _13865_ = b[423:416];
      95'b?????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13865_ = b[431:424];
      95'b????????????????????????????????????????1??????????????????????????????????????????????????????:
        _13865_ = b[439:432];
      95'b???????????????????????????????????????1???????????????????????????????????????????????????????:
        _13865_ = b[447:440];
      95'b??????????????????????????????????????1????????????????????????????????????????????????????????:
        _13865_ = b[455:448];
      95'b?????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13865_ = b[463:456];
      95'b????????????????????????????????????1??????????????????????????????????????????????????????????:
        _13865_ = b[471:464];
      95'b???????????????????????????????????1???????????????????????????????????????????????????????????:
        _13865_ = b[479:472];
      95'b??????????????????????????????????1????????????????????????????????????????????????????????????:
        _13865_ = b[487:480];
      95'b?????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13865_ = b[495:488];
      95'b????????????????????????????????1??????????????????????????????????????????????????????????????:
        _13865_ = b[503:496];
      95'b???????????????????????????????1???????????????????????????????????????????????????????????????:
        _13865_ = b[511:504];
      95'b??????????????????????????????1????????????????????????????????????????????????????????????????:
        _13865_ = b[519:512];
      95'b?????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13865_ = b[527:520];
      95'b????????????????????????????1??????????????????????????????????????????????????????????????????:
        _13865_ = b[535:528];
      95'b???????????????????????????1???????????????????????????????????????????????????????????????????:
        _13865_ = b[543:536];
      95'b??????????????????????????1????????????????????????????????????????????????????????????????????:
        _13865_ = b[551:544];
      95'b?????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13865_ = b[559:552];
      95'b????????????????????????1??????????????????????????????????????????????????????????????????????:
        _13865_ = b[567:560];
      95'b???????????????????????1???????????????????????????????????????????????????????????????????????:
        _13865_ = b[575:568];
      95'b??????????????????????1????????????????????????????????????????????????????????????????????????:
        _13865_ = b[583:576];
      95'b?????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13865_ = b[591:584];
      95'b????????????????????1??????????????????????????????????????????????????????????????????????????:
        _13865_ = b[599:592];
      95'b???????????????????1???????????????????????????????????????????????????????????????????????????:
        _13865_ = b[607:600];
      95'b??????????????????1????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[615:608];
      95'b?????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[623:616];
      95'b????????????????1??????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[631:624];
      95'b???????????????1???????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[639:632];
      95'b??????????????1????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[647:640];
      95'b?????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[655:648];
      95'b????????????1??????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[663:656];
      95'b???????????1???????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[671:664];
      95'b??????????1????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[679:672];
      95'b?????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[687:680];
      95'b????????1??????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[695:688];
      95'b???????1???????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[703:696];
      95'b??????1????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[711:704];
      95'b?????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[719:712];
      95'b????1??????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[727:720];
      95'b???1???????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[735:728];
      95'b??1????????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[743:736];
      95'b?1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[751:744];
      95'b1??????????????????????????????????????????????????????????????????????????????????????????????:
        _13865_ = b[759:752];
      default:
        _13865_ = a;
    endcase
  endfunction
  assign vec_data_094 = _13865_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744], data_d1[759:752] }, { _04536_, _04535_, _04534_, _04533_, _04532_, _04531_, _04530_, _04529_, _04528_, _04527_, _04526_, _04525_, _04524_, _04523_, _04522_, _04521_, _04520_, _04519_, _04518_, _04517_, _04516_, _04515_, _04514_, _04513_, _04512_, _04511_, _04510_, _04509_, _04508_, _04507_, _04506_, _04505_, _04504_, _04503_, _04502_, _04501_, _04500_, _04499_, _04498_, _04497_, _04496_, _04495_, _04494_, _04493_, _04492_, _04491_, _04490_, _04489_, _04488_, _04487_, _04486_, _04485_, _04484_, _04483_, _04482_, _04481_, _04480_, _04479_, _04478_, _04477_, _04476_, _04475_, _04474_, _04473_, _04472_, _04471_, _04470_, _04469_, _04468_, _04467_, _04466_, _04465_, _04464_, _04463_, _04462_, _04461_, _04460_, _04459_, _04458_, _04457_, _04456_, _04455_, _04454_, _04453_, _04452_, _04451_, _04450_, _04449_, _04448_, _04447_, _04446_, _04445_, _04444_, _04443_, _04442_ });
  assign _04442_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011111;
  assign _04443_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011110;
  assign _04444_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011101;
  assign _04445_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011100;
  assign _04446_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011011;
  assign _04447_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011010;
  assign _04448_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011001;
  assign _04449_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1011000;
  assign _04450_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010111;
  assign _04451_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010110;
  assign _04452_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010101;
  assign _04453_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010100;
  assign _04454_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010011;
  assign _04455_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010010;
  assign _04456_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010001;
  assign _04457_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1010000;
  assign _04458_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001111;
  assign _04459_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001110;
  assign _04460_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001101;
  assign _04461_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001100;
  assign _04462_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001011;
  assign _04463_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001010;
  assign _04464_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001001;
  assign _04465_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1001000;
  assign _04466_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000111;
  assign _04467_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000110;
  assign _04468_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000101;
  assign _04469_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9176|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000100;
  assign _04470_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000011;
  assign _04471_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000010;
  assign _04472_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000001;
  assign _04473_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 7'b1000000;
  assign _04474_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111111;
  assign _04475_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111110;
  assign _04476_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111101;
  assign _04477_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111100;
  assign _04478_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111011;
  assign _04479_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111010;
  assign _04480_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111001;
  assign _04481_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b111000;
  assign _04482_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110111;
  assign _04483_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110110;
  assign _04484_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110101;
  assign _04485_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110100;
  assign _04486_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110011;
  assign _04487_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110010;
  assign _04488_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110001;
  assign _04489_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b110000;
  assign _04490_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101111;
  assign _04491_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101110;
  assign _04492_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101101;
  assign _04493_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101100;
  assign _04494_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101011;
  assign _04495_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101010;
  assign _04496_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101001;
  assign _04497_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b101000;
  assign _04498_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100111;
  assign _04499_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100110;
  assign _04500_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100101;
  assign _04501_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100100;
  assign _04502_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100011;
  assign _04503_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100010;
  assign _04504_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100001;
  assign _04505_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 6'b100000;
  assign _04506_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11111;
  assign _04507_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11110;
  assign _04508_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11101;
  assign _04509_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11100;
  assign _04510_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11011;
  assign _04511_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11010;
  assign _04512_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11001;
  assign _04513_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b11000;
  assign _04514_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10111;
  assign _04515_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10110;
  assign _04516_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10101;
  assign _04517_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10100;
  assign _04518_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10011;
  assign _04519_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10010;
  assign _04520_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10001;
  assign _04521_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 5'b10000;
  assign _04522_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1111;
  assign _04523_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1110;
  assign _04524_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1101;
  assign _04525_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1100;
  assign _04526_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1011;
  assign _04527_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1010;
  assign _04528_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1001;
  assign _04529_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 4'b1000;
  assign _04530_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 3'b111;
  assign _04531_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 3'b110;
  assign _04532_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 3'b101;
  assign _04533_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 3'b100;
  assign _04534_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 2'b11;
  assign _04535_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 2'b10;
  assign _04536_ = vec_sum_094_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9108" *) 1'b1;
  function [7:0] _13961_;
    input [7:0] a;
    input [751:0] b;
    input [93:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *)
    (* parallel_case *)
    casez (s)
      94'b?????????????????????????????????????????????????????????????????????????????????????????????1:
        _13961_ = b[7:0];
      94'b????????????????????????????????????????????????????????????????????????????????????????????1?:
        _13961_ = b[15:8];
      94'b???????????????????????????????????????????????????????????????????????????????????????????1??:
        _13961_ = b[23:16];
      94'b??????????????????????????????????????????????????????????????????????????????????????????1???:
        _13961_ = b[31:24];
      94'b?????????????????????????????????????????????????????????????????????????????????????????1????:
        _13961_ = b[39:32];
      94'b????????????????????????????????????????????????????????????????????????????????????????1?????:
        _13961_ = b[47:40];
      94'b???????????????????????????????????????????????????????????????????????????????????????1??????:
        _13961_ = b[55:48];
      94'b??????????????????????????????????????????????????????????????????????????????????????1???????:
        _13961_ = b[63:56];
      94'b?????????????????????????????????????????????????????????????????????????????????????1????????:
        _13961_ = b[71:64];
      94'b????????????????????????????????????????????????????????????????????????????????????1?????????:
        _13961_ = b[79:72];
      94'b???????????????????????????????????????????????????????????????????????????????????1??????????:
        _13961_ = b[87:80];
      94'b??????????????????????????????????????????????????????????????????????????????????1???????????:
        _13961_ = b[95:88];
      94'b?????????????????????????????????????????????????????????????????????????????????1????????????:
        _13961_ = b[103:96];
      94'b????????????????????????????????????????????????????????????????????????????????1?????????????:
        _13961_ = b[111:104];
      94'b???????????????????????????????????????????????????????????????????????????????1??????????????:
        _13961_ = b[119:112];
      94'b??????????????????????????????????????????????????????????????????????????????1???????????????:
        _13961_ = b[127:120];
      94'b?????????????????????????????????????????????????????????????????????????????1????????????????:
        _13961_ = b[135:128];
      94'b????????????????????????????????????????????????????????????????????????????1?????????????????:
        _13961_ = b[143:136];
      94'b???????????????????????????????????????????????????????????????????????????1??????????????????:
        _13961_ = b[151:144];
      94'b??????????????????????????????????????????????????????????????????????????1???????????????????:
        _13961_ = b[159:152];
      94'b?????????????????????????????????????????????????????????????????????????1????????????????????:
        _13961_ = b[167:160];
      94'b????????????????????????????????????????????????????????????????????????1?????????????????????:
        _13961_ = b[175:168];
      94'b???????????????????????????????????????????????????????????????????????1??????????????????????:
        _13961_ = b[183:176];
      94'b??????????????????????????????????????????????????????????????????????1???????????????????????:
        _13961_ = b[191:184];
      94'b?????????????????????????????????????????????????????????????????????1????????????????????????:
        _13961_ = b[199:192];
      94'b????????????????????????????????????????????????????????????????????1?????????????????????????:
        _13961_ = b[207:200];
      94'b???????????????????????????????????????????????????????????????????1??????????????????????????:
        _13961_ = b[215:208];
      94'b??????????????????????????????????????????????????????????????????1???????????????????????????:
        _13961_ = b[223:216];
      94'b?????????????????????????????????????????????????????????????????1????????????????????????????:
        _13961_ = b[231:224];
      94'b????????????????????????????????????????????????????????????????1?????????????????????????????:
        _13961_ = b[239:232];
      94'b???????????????????????????????????????????????????????????????1??????????????????????????????:
        _13961_ = b[247:240];
      94'b??????????????????????????????????????????????????????????????1???????????????????????????????:
        _13961_ = b[255:248];
      94'b?????????????????????????????????????????????????????????????1????????????????????????????????:
        _13961_ = b[263:256];
      94'b????????????????????????????????????????????????????????????1?????????????????????????????????:
        _13961_ = b[271:264];
      94'b???????????????????????????????????????????????????????????1??????????????????????????????????:
        _13961_ = b[279:272];
      94'b??????????????????????????????????????????????????????????1???????????????????????????????????:
        _13961_ = b[287:280];
      94'b?????????????????????????????????????????????????????????1????????????????????????????????????:
        _13961_ = b[295:288];
      94'b????????????????????????????????????????????????????????1?????????????????????????????????????:
        _13961_ = b[303:296];
      94'b???????????????????????????????????????????????????????1??????????????????????????????????????:
        _13961_ = b[311:304];
      94'b??????????????????????????????????????????????????????1???????????????????????????????????????:
        _13961_ = b[319:312];
      94'b?????????????????????????????????????????????????????1????????????????????????????????????????:
        _13961_ = b[327:320];
      94'b????????????????????????????????????????????????????1?????????????????????????????????????????:
        _13961_ = b[335:328];
      94'b???????????????????????????????????????????????????1??????????????????????????????????????????:
        _13961_ = b[343:336];
      94'b??????????????????????????????????????????????????1???????????????????????????????????????????:
        _13961_ = b[351:344];
      94'b?????????????????????????????????????????????????1????????????????????????????????????????????:
        _13961_ = b[359:352];
      94'b????????????????????????????????????????????????1?????????????????????????????????????????????:
        _13961_ = b[367:360];
      94'b???????????????????????????????????????????????1??????????????????????????????????????????????:
        _13961_ = b[375:368];
      94'b??????????????????????????????????????????????1???????????????????????????????????????????????:
        _13961_ = b[383:376];
      94'b?????????????????????????????????????????????1????????????????????????????????????????????????:
        _13961_ = b[391:384];
      94'b????????????????????????????????????????????1?????????????????????????????????????????????????:
        _13961_ = b[399:392];
      94'b???????????????????????????????????????????1??????????????????????????????????????????????????:
        _13961_ = b[407:400];
      94'b??????????????????????????????????????????1???????????????????????????????????????????????????:
        _13961_ = b[415:408];
      94'b?????????????????????????????????????????1????????????????????????????????????????????????????:
        _13961_ = b[423:416];
      94'b????????????????????????????????????????1?????????????????????????????????????????????????????:
        _13961_ = b[431:424];
      94'b???????????????????????????????????????1??????????????????????????????????????????????????????:
        _13961_ = b[439:432];
      94'b??????????????????????????????????????1???????????????????????????????????????????????????????:
        _13961_ = b[447:440];
      94'b?????????????????????????????????????1????????????????????????????????????????????????????????:
        _13961_ = b[455:448];
      94'b????????????????????????????????????1?????????????????????????????????????????????????????????:
        _13961_ = b[463:456];
      94'b???????????????????????????????????1??????????????????????????????????????????????????????????:
        _13961_ = b[471:464];
      94'b??????????????????????????????????1???????????????????????????????????????????????????????????:
        _13961_ = b[479:472];
      94'b?????????????????????????????????1????????????????????????????????????????????????????????????:
        _13961_ = b[487:480];
      94'b????????????????????????????????1?????????????????????????????????????????????????????????????:
        _13961_ = b[495:488];
      94'b???????????????????????????????1??????????????????????????????????????????????????????????????:
        _13961_ = b[503:496];
      94'b??????????????????????????????1???????????????????????????????????????????????????????????????:
        _13961_ = b[511:504];
      94'b?????????????????????????????1????????????????????????????????????????????????????????????????:
        _13961_ = b[519:512];
      94'b????????????????????????????1?????????????????????????????????????????????????????????????????:
        _13961_ = b[527:520];
      94'b???????????????????????????1??????????????????????????????????????????????????????????????????:
        _13961_ = b[535:528];
      94'b??????????????????????????1???????????????????????????????????????????????????????????????????:
        _13961_ = b[543:536];
      94'b?????????????????????????1????????????????????????????????????????????????????????????????????:
        _13961_ = b[551:544];
      94'b????????????????????????1?????????????????????????????????????????????????????????????????????:
        _13961_ = b[559:552];
      94'b???????????????????????1??????????????????????????????????????????????????????????????????????:
        _13961_ = b[567:560];
      94'b??????????????????????1???????????????????????????????????????????????????????????????????????:
        _13961_ = b[575:568];
      94'b?????????????????????1????????????????????????????????????????????????????????????????????????:
        _13961_ = b[583:576];
      94'b????????????????????1?????????????????????????????????????????????????????????????????????????:
        _13961_ = b[591:584];
      94'b???????????????????1??????????????????????????????????????????????????????????????????????????:
        _13961_ = b[599:592];
      94'b??????????????????1???????????????????????????????????????????????????????????????????????????:
        _13961_ = b[607:600];
      94'b?????????????????1????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[615:608];
      94'b????????????????1?????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[623:616];
      94'b???????????????1??????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[631:624];
      94'b??????????????1???????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[639:632];
      94'b?????????????1????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[647:640];
      94'b????????????1?????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[655:648];
      94'b???????????1??????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[663:656];
      94'b??????????1???????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[671:664];
      94'b?????????1????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[679:672];
      94'b????????1?????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[687:680];
      94'b???????1??????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[695:688];
      94'b??????1???????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[703:696];
      94'b?????1????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[711:704];
      94'b????1?????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[719:712];
      94'b???1??????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[727:720];
      94'b??1???????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[735:728];
      94'b?1????????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[743:736];
      94'b1?????????????????????????????????????????????????????????????????????????????????????????????:
        _13961_ = b[751:744];
      default:
        _13961_ = a;
    endcase
  endfunction
  assign vec_data_093 = _13961_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736], data_d1[751:744] }, { _04630_, _04629_, _04628_, _04627_, _04626_, _04625_, _04624_, _04623_, _04622_, _04621_, _04620_, _04619_, _04618_, _04617_, _04616_, _04615_, _04614_, _04613_, _04612_, _04611_, _04610_, _04609_, _04608_, _04607_, _04606_, _04605_, _04604_, _04603_, _04602_, _04601_, _04600_, _04599_, _04598_, _04597_, _04596_, _04595_, _04594_, _04593_, _04592_, _04591_, _04590_, _04589_, _04588_, _04587_, _04586_, _04585_, _04584_, _04583_, _04582_, _04581_, _04580_, _04579_, _04578_, _04577_, _04576_, _04575_, _04574_, _04573_, _04572_, _04571_, _04570_, _04569_, _04568_, _04567_, _04566_, _04565_, _04564_, _04563_, _04562_, _04561_, _04560_, _04559_, _04558_, _04557_, _04556_, _04555_, _04554_, _04553_, _04552_, _04551_, _04550_, _04549_, _04548_, _04547_, _04546_, _04545_, _04544_, _04543_, _04542_, _04541_, _04540_, _04539_, _04538_, _04537_ });
  assign _04537_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011110;
  assign _04538_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011101;
  assign _04539_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011100;
  assign _04540_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011011;
  assign _04541_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011010;
  assign _04542_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011001;
  assign _04543_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1011000;
  assign _04544_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010111;
  assign _04545_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010110;
  assign _04546_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010101;
  assign _04547_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010100;
  assign _04548_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010011;
  assign _04549_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010010;
  assign _04550_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010001;
  assign _04551_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1010000;
  assign _04552_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001111;
  assign _04553_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001110;
  assign _04554_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001101;
  assign _04555_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001100;
  assign _04556_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001011;
  assign _04557_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001010;
  assign _04558_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001001;
  assign _04559_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1001000;
  assign _04560_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000111;
  assign _04561_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000110;
  assign _04562_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000101;
  assign _04563_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000100;
  assign _04564_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000011;
  assign _04565_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000010;
  assign _04566_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000001;
  assign _04567_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 7'b1000000;
  assign _04568_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111111;
  assign _04569_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111110;
  assign _04570_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111101;
  assign _04571_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111100;
  assign _04572_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111011;
  assign _04573_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111010;
  assign _04574_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111001;
  assign _04575_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b111000;
  assign _04576_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110111;
  assign _04577_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110110;
  assign _04578_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110101;
  assign _04579_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110100;
  assign _04580_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110011;
  assign _04581_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110010;
  assign _04582_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110001;
  assign _04583_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b110000;
  assign _04584_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101111;
  assign _04585_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101110;
  assign _04586_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101101;
  assign _04587_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101100;
  assign _04588_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101011;
  assign _04589_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101010;
  assign _04590_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101001;
  assign _04591_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b101000;
  assign _04592_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100111;
  assign _04593_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100110;
  assign _04594_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100101;
  assign _04595_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100100;
  assign _04596_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100011;
  assign _04597_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100010;
  assign _04598_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100001;
  assign _04599_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 6'b100000;
  assign _04600_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11111;
  assign _04601_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11110;
  assign _04602_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11101;
  assign _04603_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11100;
  assign _04604_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11011;
  assign _04605_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11010;
  assign _04606_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11001;
  assign _04607_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b11000;
  assign _04608_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10111;
  assign _04609_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10110;
  assign _04610_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10101;
  assign _04611_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10100;
  assign _04612_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10011;
  assign _04613_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10010;
  assign _04614_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10001;
  assign _04615_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 5'b10000;
  assign _04616_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1111;
  assign _04617_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1110;
  assign _04618_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1101;
  assign _04619_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1100;
  assign _04620_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1011;
  assign _04621_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1010;
  assign _04622_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1001;
  assign _04623_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 4'b1000;
  assign _04624_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 3'b111;
  assign _04625_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 3'b110;
  assign _04626_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 3'b101;
  assign _04627_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 3'b100;
  assign _04628_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 2'b11;
  assign _04629_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 2'b10;
  assign _04630_ = vec_sum_093_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:9006" *) 1'b1;
  function [7:0] _14056_;
    input [7:0] a;
    input [743:0] b;
    input [92:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *)
    (* parallel_case *)
    casez (s)
      93'b????????????????????????????????????????????????????????????????????????????????????????????1:
        _14056_ = b[7:0];
      93'b???????????????????????????????????????????????????????????????????????????????????????????1?:
        _14056_ = b[15:8];
      93'b??????????????????????????????????????????????????????????????????????????????????????????1??:
        _14056_ = b[23:16];
      93'b?????????????????????????????????????????????????????????????????????????????????????????1???:
        _14056_ = b[31:24];
      93'b????????????????????????????????????????????????????????????????????????????????????????1????:
        _14056_ = b[39:32];
      93'b???????????????????????????????????????????????????????????????????????????????????????1?????:
        _14056_ = b[47:40];
      93'b??????????????????????????????????????????????????????????????????????????????????????1??????:
        _14056_ = b[55:48];
      93'b?????????????????????????????????????????????????????????????????????????????????????1???????:
        _14056_ = b[63:56];
      93'b????????????????????????????????????????????????????????????????????????????????????1????????:
        _14056_ = b[71:64];
      93'b???????????????????????????????????????????????????????????????????????????????????1?????????:
        _14056_ = b[79:72];
      93'b??????????????????????????????????????????????????????????????????????????????????1??????????:
        _14056_ = b[87:80];
      93'b?????????????????????????????????????????????????????????????????????????????????1???????????:
        _14056_ = b[95:88];
      93'b????????????????????????????????????????????????????????????????????????????????1????????????:
        _14056_ = b[103:96];
      93'b???????????????????????????????????????????????????????????????????????????????1?????????????:
        _14056_ = b[111:104];
      93'b??????????????????????????????????????????????????????????????????????????????1??????????????:
        _14056_ = b[119:112];
      93'b?????????????????????????????????????????????????????????????????????????????1???????????????:
        _14056_ = b[127:120];
      93'b????????????????????????????????????????????????????????????????????????????1????????????????:
        _14056_ = b[135:128];
      93'b???????????????????????????????????????????????????????????????????????????1?????????????????:
        _14056_ = b[143:136];
      93'b??????????????????????????????????????????????????????????????????????????1??????????????????:
        _14056_ = b[151:144];
      93'b?????????????????????????????????????????????????????????????????????????1???????????????????:
        _14056_ = b[159:152];
      93'b????????????????????????????????????????????????????????????????????????1????????????????????:
        _14056_ = b[167:160];
      93'b???????????????????????????????????????????????????????????????????????1?????????????????????:
        _14056_ = b[175:168];
      93'b??????????????????????????????????????????????????????????????????????1??????????????????????:
        _14056_ = b[183:176];
      93'b?????????????????????????????????????????????????????????????????????1???????????????????????:
        _14056_ = b[191:184];
      93'b????????????????????????????????????????????????????????????????????1????????????????????????:
        _14056_ = b[199:192];
      93'b???????????????????????????????????????????????????????????????????1?????????????????????????:
        _14056_ = b[207:200];
      93'b??????????????????????????????????????????????????????????????????1??????????????????????????:
        _14056_ = b[215:208];
      93'b?????????????????????????????????????????????????????????????????1???????????????????????????:
        _14056_ = b[223:216];
      93'b????????????????????????????????????????????????????????????????1????????????????????????????:
        _14056_ = b[231:224];
      93'b???????????????????????????????????????????????????????????????1?????????????????????????????:
        _14056_ = b[239:232];
      93'b??????????????????????????????????????????????????????????????1??????????????????????????????:
        _14056_ = b[247:240];
      93'b?????????????????????????????????????????????????????????????1???????????????????????????????:
        _14056_ = b[255:248];
      93'b????????????????????????????????????????????????????????????1????????????????????????????????:
        _14056_ = b[263:256];
      93'b???????????????????????????????????????????????????????????1?????????????????????????????????:
        _14056_ = b[271:264];
      93'b??????????????????????????????????????????????????????????1??????????????????????????????????:
        _14056_ = b[279:272];
      93'b?????????????????????????????????????????????????????????1???????????????????????????????????:
        _14056_ = b[287:280];
      93'b????????????????????????????????????????????????????????1????????????????????????????????????:
        _14056_ = b[295:288];
      93'b???????????????????????????????????????????????????????1?????????????????????????????????????:
        _14056_ = b[303:296];
      93'b??????????????????????????????????????????????????????1??????????????????????????????????????:
        _14056_ = b[311:304];
      93'b?????????????????????????????????????????????????????1???????????????????????????????????????:
        _14056_ = b[319:312];
      93'b????????????????????????????????????????????????????1????????????????????????????????????????:
        _14056_ = b[327:320];
      93'b???????????????????????????????????????????????????1?????????????????????????????????????????:
        _14056_ = b[335:328];
      93'b??????????????????????????????????????????????????1??????????????????????????????????????????:
        _14056_ = b[343:336];
      93'b?????????????????????????????????????????????????1???????????????????????????????????????????:
        _14056_ = b[351:344];
      93'b????????????????????????????????????????????????1????????????????????????????????????????????:
        _14056_ = b[359:352];
      93'b???????????????????????????????????????????????1?????????????????????????????????????????????:
        _14056_ = b[367:360];
      93'b??????????????????????????????????????????????1??????????????????????????????????????????????:
        _14056_ = b[375:368];
      93'b?????????????????????????????????????????????1???????????????????????????????????????????????:
        _14056_ = b[383:376];
      93'b????????????????????????????????????????????1????????????????????????????????????????????????:
        _14056_ = b[391:384];
      93'b???????????????????????????????????????????1?????????????????????????????????????????????????:
        _14056_ = b[399:392];
      93'b??????????????????????????????????????????1??????????????????????????????????????????????????:
        _14056_ = b[407:400];
      93'b?????????????????????????????????????????1???????????????????????????????????????????????????:
        _14056_ = b[415:408];
      93'b????????????????????????????????????????1????????????????????????????????????????????????????:
        _14056_ = b[423:416];
      93'b???????????????????????????????????????1?????????????????????????????????????????????????????:
        _14056_ = b[431:424];
      93'b??????????????????????????????????????1??????????????????????????????????????????????????????:
        _14056_ = b[439:432];
      93'b?????????????????????????????????????1???????????????????????????????????????????????????????:
        _14056_ = b[447:440];
      93'b????????????????????????????????????1????????????????????????????????????????????????????????:
        _14056_ = b[455:448];
      93'b???????????????????????????????????1?????????????????????????????????????????????????????????:
        _14056_ = b[463:456];
      93'b??????????????????????????????????1??????????????????????????????????????????????????????????:
        _14056_ = b[471:464];
      93'b?????????????????????????????????1???????????????????????????????????????????????????????????:
        _14056_ = b[479:472];
      93'b????????????????????????????????1????????????????????????????????????????????????????????????:
        _14056_ = b[487:480];
      93'b???????????????????????????????1?????????????????????????????????????????????????????????????:
        _14056_ = b[495:488];
      93'b??????????????????????????????1??????????????????????????????????????????????????????????????:
        _14056_ = b[503:496];
      93'b?????????????????????????????1???????????????????????????????????????????????????????????????:
        _14056_ = b[511:504];
      93'b????????????????????????????1????????????????????????????????????????????????????????????????:
        _14056_ = b[519:512];
      93'b???????????????????????????1?????????????????????????????????????????????????????????????????:
        _14056_ = b[527:520];
      93'b??????????????????????????1??????????????????????????????????????????????????????????????????:
        _14056_ = b[535:528];
      93'b?????????????????????????1???????????????????????????????????????????????????????????????????:
        _14056_ = b[543:536];
      93'b????????????????????????1????????????????????????????????????????????????????????????????????:
        _14056_ = b[551:544];
      93'b???????????????????????1?????????????????????????????????????????????????????????????????????:
        _14056_ = b[559:552];
      93'b??????????????????????1??????????????????????????????????????????????????????????????????????:
        _14056_ = b[567:560];
      93'b?????????????????????1???????????????????????????????????????????????????????????????????????:
        _14056_ = b[575:568];
      93'b????????????????????1????????????????????????????????????????????????????????????????????????:
        _14056_ = b[583:576];
      93'b???????????????????1?????????????????????????????????????????????????????????????????????????:
        _14056_ = b[591:584];
      93'b??????????????????1??????????????????????????????????????????????????????????????????????????:
        _14056_ = b[599:592];
      93'b?????????????????1???????????????????????????????????????????????????????????????????????????:
        _14056_ = b[607:600];
      93'b????????????????1????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[615:608];
      93'b???????????????1?????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[623:616];
      93'b??????????????1??????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[631:624];
      93'b?????????????1???????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[639:632];
      93'b????????????1????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[647:640];
      93'b???????????1?????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[655:648];
      93'b??????????1??????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[663:656];
      93'b?????????1???????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[671:664];
      93'b????????1????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[679:672];
      93'b???????1?????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[687:680];
      93'b??????1??????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[695:688];
      93'b?????1???????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[703:696];
      93'b????1????????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[711:704];
      93'b???1?????????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[719:712];
      93'b??1??????????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[727:720];
      93'b?1???????????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[735:728];
      93'b1????????????????????????????????????????????????????????????????????????????????????????????:
        _14056_ = b[743:736];
      default:
        _14056_ = a;
    endcase
  endfunction
  assign vec_data_092 = _14056_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728], data_d1[743:736] }, { _04723_, _04722_, _04721_, _04720_, _04719_, _04718_, _04717_, _04716_, _04715_, _04714_, _04713_, _04712_, _04711_, _04710_, _04709_, _04708_, _04707_, _04706_, _04705_, _04704_, _04703_, _04702_, _04701_, _04700_, _04699_, _04698_, _04697_, _04696_, _04695_, _04694_, _04693_, _04692_, _04691_, _04690_, _04689_, _04688_, _04687_, _04686_, _04685_, _04684_, _04683_, _04682_, _04681_, _04680_, _04679_, _04678_, _04677_, _04676_, _04675_, _04674_, _04673_, _04672_, _04671_, _04670_, _04669_, _04668_, _04667_, _04666_, _04665_, _04664_, _04663_, _04662_, _04661_, _04660_, _04659_, _04658_, _04657_, _04656_, _04655_, _04654_, _04653_, _04652_, _04651_, _04650_, _04649_, _04648_, _04647_, _04646_, _04645_, _04644_, _04643_, _04642_, _04641_, _04640_, _04639_, _04638_, _04637_, _04636_, _04635_, _04634_, _04633_, _04632_, _04631_ });
  assign _04631_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011101;
  assign _04632_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011100;
  assign _04633_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011011;
  assign _04634_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011010;
  assign _04635_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011001;
  assign _04636_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1011000;
  assign _04637_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010111;
  assign _04638_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010110;
  assign _04639_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010101;
  assign _04640_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010100;
  assign _04641_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010011;
  assign _04642_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010010;
  assign _04643_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010001;
  assign _04644_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1010000;
  assign _04645_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001111;
  assign _04646_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001110;
  assign _04647_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001101;
  assign _04648_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001100;
  assign _04649_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001011;
  assign _04650_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001010;
  assign _04651_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001001;
  assign _04652_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1001000;
  assign _04653_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000111;
  assign _04654_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000110;
  assign _04655_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000101;
  assign _04656_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000100;
  assign _04657_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000011;
  assign _04658_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000010;
  assign _04659_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000001;
  assign _04660_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 7'b1000000;
  assign _04661_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111111;
  assign _04662_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111110;
  assign _04663_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111101;
  assign _04664_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111100;
  assign _04665_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111011;
  assign _04666_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111010;
  assign _04667_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111001;
  assign _04668_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b111000;
  assign _04669_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110111;
  assign _04670_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110110;
  assign _04671_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110101;
  assign _04672_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110100;
  assign _04673_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110011;
  assign _04674_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110010;
  assign _04675_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110001;
  assign _04676_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b110000;
  assign _04677_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101111;
  assign _04678_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101110;
  assign _04679_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101101;
  assign _04680_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101100;
  assign _04681_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101011;
  assign _04682_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101010;
  assign _04683_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101001;
  assign _04684_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b101000;
  assign _04685_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100111;
  assign _04686_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100110;
  assign _04687_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100101;
  assign _04688_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100100;
  assign _04689_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100011;
  assign _04690_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100010;
  assign _04691_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100001;
  assign _04692_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 6'b100000;
  assign _04693_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11111;
  assign _04694_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11110;
  assign _04695_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11101;
  assign _04696_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11100;
  assign _04697_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11011;
  assign _04698_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11010;
  assign _04699_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11001;
  assign _04700_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b11000;
  assign _04701_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10111;
  assign _04702_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10110;
  assign _04703_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10101;
  assign _04704_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10100;
  assign _04705_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10011;
  assign _04706_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10010;
  assign _04707_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10001;
  assign _04708_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 5'b10000;
  assign _04709_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1111;
  assign _04710_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1110;
  assign _04711_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1101;
  assign _04712_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1100;
  assign _04713_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1011;
  assign _04714_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1010;
  assign _04715_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1001;
  assign _04716_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 4'b1000;
  assign _04717_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 3'b111;
  assign _04718_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 3'b110;
  assign _04719_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 3'b101;
  assign _04720_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 3'b100;
  assign _04721_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 2'b11;
  assign _04722_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 2'b10;
  assign _04723_ = vec_sum_092_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8905" *) 1'b1;
  function [7:0] _14150_;
    input [7:0] a;
    input [735:0] b;
    input [91:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *)
    (* parallel_case *)
    casez (s)
      92'b???????????????????????????????????????????????????????????????????????????????????????????1:
        _14150_ = b[7:0];
      92'b??????????????????????????????????????????????????????????????????????????????????????????1?:
        _14150_ = b[15:8];
      92'b?????????????????????????????????????????????????????????????????????????????????????????1??:
        _14150_ = b[23:16];
      92'b????????????????????????????????????????????????????????????????????????????????????????1???:
        _14150_ = b[31:24];
      92'b???????????????????????????????????????????????????????????????????????????????????????1????:
        _14150_ = b[39:32];
      92'b??????????????????????????????????????????????????????????????????????????????????????1?????:
        _14150_ = b[47:40];
      92'b?????????????????????????????????????????????????????????????????????????????????????1??????:
        _14150_ = b[55:48];
      92'b????????????????????????????????????????????????????????????????????????????????????1???????:
        _14150_ = b[63:56];
      92'b???????????????????????????????????????????????????????????????????????????????????1????????:
        _14150_ = b[71:64];
      92'b??????????????????????????????????????????????????????????????????????????????????1?????????:
        _14150_ = b[79:72];
      92'b?????????????????????????????????????????????????????????????????????????????????1??????????:
        _14150_ = b[87:80];
      92'b????????????????????????????????????????????????????????????????????????????????1???????????:
        _14150_ = b[95:88];
      92'b???????????????????????????????????????????????????????????????????????????????1????????????:
        _14150_ = b[103:96];
      92'b??????????????????????????????????????????????????????????????????????????????1?????????????:
        _14150_ = b[111:104];
      92'b?????????????????????????????????????????????????????????????????????????????1??????????????:
        _14150_ = b[119:112];
      92'b????????????????????????????????????????????????????????????????????????????1???????????????:
        _14150_ = b[127:120];
      92'b???????????????????????????????????????????????????????????????????????????1????????????????:
        _14150_ = b[135:128];
      92'b??????????????????????????????????????????????????????????????????????????1?????????????????:
        _14150_ = b[143:136];
      92'b?????????????????????????????????????????????????????????????????????????1??????????????????:
        _14150_ = b[151:144];
      92'b????????????????????????????????????????????????????????????????????????1???????????????????:
        _14150_ = b[159:152];
      92'b???????????????????????????????????????????????????????????????????????1????????????????????:
        _14150_ = b[167:160];
      92'b??????????????????????????????????????????????????????????????????????1?????????????????????:
        _14150_ = b[175:168];
      92'b?????????????????????????????????????????????????????????????????????1??????????????????????:
        _14150_ = b[183:176];
      92'b????????????????????????????????????????????????????????????????????1???????????????????????:
        _14150_ = b[191:184];
      92'b???????????????????????????????????????????????????????????????????1????????????????????????:
        _14150_ = b[199:192];
      92'b??????????????????????????????????????????????????????????????????1?????????????????????????:
        _14150_ = b[207:200];
      92'b?????????????????????????????????????????????????????????????????1??????????????????????????:
        _14150_ = b[215:208];
      92'b????????????????????????????????????????????????????????????????1???????????????????????????:
        _14150_ = b[223:216];
      92'b???????????????????????????????????????????????????????????????1????????????????????????????:
        _14150_ = b[231:224];
      92'b??????????????????????????????????????????????????????????????1?????????????????????????????:
        _14150_ = b[239:232];
      92'b?????????????????????????????????????????????????????????????1??????????????????????????????:
        _14150_ = b[247:240];
      92'b????????????????????????????????????????????????????????????1???????????????????????????????:
        _14150_ = b[255:248];
      92'b???????????????????????????????????????????????????????????1????????????????????????????????:
        _14150_ = b[263:256];
      92'b??????????????????????????????????????????????????????????1?????????????????????????????????:
        _14150_ = b[271:264];
      92'b?????????????????????????????????????????????????????????1??????????????????????????????????:
        _14150_ = b[279:272];
      92'b????????????????????????????????????????????????????????1???????????????????????????????????:
        _14150_ = b[287:280];
      92'b???????????????????????????????????????????????????????1????????????????????????????????????:
        _14150_ = b[295:288];
      92'b??????????????????????????????????????????????????????1?????????????????????????????????????:
        _14150_ = b[303:296];
      92'b?????????????????????????????????????????????????????1??????????????????????????????????????:
        _14150_ = b[311:304];
      92'b????????????????????????????????????????????????????1???????????????????????????????????????:
        _14150_ = b[319:312];
      92'b???????????????????????????????????????????????????1????????????????????????????????????????:
        _14150_ = b[327:320];
      92'b??????????????????????????????????????????????????1?????????????????????????????????????????:
        _14150_ = b[335:328];
      92'b?????????????????????????????????????????????????1??????????????????????????????????????????:
        _14150_ = b[343:336];
      92'b????????????????????????????????????????????????1???????????????????????????????????????????:
        _14150_ = b[351:344];
      92'b???????????????????????????????????????????????1????????????????????????????????????????????:
        _14150_ = b[359:352];
      92'b??????????????????????????????????????????????1?????????????????????????????????????????????:
        _14150_ = b[367:360];
      92'b?????????????????????????????????????????????1??????????????????????????????????????????????:
        _14150_ = b[375:368];
      92'b????????????????????????????????????????????1???????????????????????????????????????????????:
        _14150_ = b[383:376];
      92'b???????????????????????????????????????????1????????????????????????????????????????????????:
        _14150_ = b[391:384];
      92'b??????????????????????????????????????????1?????????????????????????????????????????????????:
        _14150_ = b[399:392];
      92'b?????????????????????????????????????????1??????????????????????????????????????????????????:
        _14150_ = b[407:400];
      92'b????????????????????????????????????????1???????????????????????????????????????????????????:
        _14150_ = b[415:408];
      92'b???????????????????????????????????????1????????????????????????????????????????????????????:
        _14150_ = b[423:416];
      92'b??????????????????????????????????????1?????????????????????????????????????????????????????:
        _14150_ = b[431:424];
      92'b?????????????????????????????????????1??????????????????????????????????????????????????????:
        _14150_ = b[439:432];
      92'b????????????????????????????????????1???????????????????????????????????????????????????????:
        _14150_ = b[447:440];
      92'b???????????????????????????????????1????????????????????????????????????????????????????????:
        _14150_ = b[455:448];
      92'b??????????????????????????????????1?????????????????????????????????????????????????????????:
        _14150_ = b[463:456];
      92'b?????????????????????????????????1??????????????????????????????????????????????????????????:
        _14150_ = b[471:464];
      92'b????????????????????????????????1???????????????????????????????????????????????????????????:
        _14150_ = b[479:472];
      92'b???????????????????????????????1????????????????????????????????????????????????????????????:
        _14150_ = b[487:480];
      92'b??????????????????????????????1?????????????????????????????????????????????????????????????:
        _14150_ = b[495:488];
      92'b?????????????????????????????1??????????????????????????????????????????????????????????????:
        _14150_ = b[503:496];
      92'b????????????????????????????1???????????????????????????????????????????????????????????????:
        _14150_ = b[511:504];
      92'b???????????????????????????1????????????????????????????????????????????????????????????????:
        _14150_ = b[519:512];
      92'b??????????????????????????1?????????????????????????????????????????????????????????????????:
        _14150_ = b[527:520];
      92'b?????????????????????????1??????????????????????????????????????????????????????????????????:
        _14150_ = b[535:528];
      92'b????????????????????????1???????????????????????????????????????????????????????????????????:
        _14150_ = b[543:536];
      92'b???????????????????????1????????????????????????????????????????????????????????????????????:
        _14150_ = b[551:544];
      92'b??????????????????????1?????????????????????????????????????????????????????????????????????:
        _14150_ = b[559:552];
      92'b?????????????????????1??????????????????????????????????????????????????????????????????????:
        _14150_ = b[567:560];
      92'b????????????????????1???????????????????????????????????????????????????????????????????????:
        _14150_ = b[575:568];
      92'b???????????????????1????????????????????????????????????????????????????????????????????????:
        _14150_ = b[583:576];
      92'b??????????????????1?????????????????????????????????????????????????????????????????????????:
        _14150_ = b[591:584];
      92'b?????????????????1??????????????????????????????????????????????????????????????????????????:
        _14150_ = b[599:592];
      92'b????????????????1???????????????????????????????????????????????????????????????????????????:
        _14150_ = b[607:600];
      92'b???????????????1????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[615:608];
      92'b??????????????1?????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[623:616];
      92'b?????????????1??????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[631:624];
      92'b????????????1???????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[639:632];
      92'b???????????1????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[647:640];
      92'b??????????1?????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[655:648];
      92'b?????????1??????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[663:656];
      92'b????????1???????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[671:664];
      92'b???????1????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[679:672];
      92'b??????1?????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[687:680];
      92'b?????1??????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[695:688];
      92'b????1???????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[703:696];
      92'b???1????????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[711:704];
      92'b??1?????????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[719:712];
      92'b?1??????????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[727:720];
      92'b1???????????????????????????????????????????????????????????????????????????????????????????:
        _14150_ = b[735:728];
      default:
        _14150_ = a;
    endcase
  endfunction
  assign vec_data_091 = _14150_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720], data_d1[735:728] }, { _04815_, _04814_, _04813_, _04812_, _04811_, _04810_, _04809_, _04808_, _04807_, _04806_, _04805_, _04804_, _04803_, _04802_, _04801_, _04800_, _04799_, _04798_, _04797_, _04796_, _04795_, _04794_, _04793_, _04792_, _04791_, _04790_, _04789_, _04788_, _04787_, _04786_, _04785_, _04784_, _04783_, _04782_, _04781_, _04780_, _04779_, _04778_, _04777_, _04776_, _04775_, _04774_, _04773_, _04772_, _04771_, _04770_, _04769_, _04768_, _04767_, _04766_, _04765_, _04764_, _04763_, _04762_, _04761_, _04760_, _04759_, _04758_, _04757_, _04756_, _04755_, _04754_, _04753_, _04752_, _04751_, _04750_, _04749_, _04748_, _04747_, _04746_, _04745_, _04744_, _04743_, _04742_, _04741_, _04740_, _04739_, _04738_, _04737_, _04736_, _04735_, _04734_, _04733_, _04732_, _04731_, _04730_, _04729_, _04728_, _04727_, _04726_, _04725_, _04724_ });
  assign _04724_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1011100;
  assign _04725_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1011011;
  assign _04726_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1011010;
  assign _04727_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1011001;
  assign _04728_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1011000;
  assign _04729_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010111;
  assign _04730_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010110;
  assign _04731_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010101;
  assign _04732_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010100;
  assign _04733_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010011;
  assign _04734_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010010;
  assign _04735_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010001;
  assign _04736_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1010000;
  assign _04737_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001111;
  assign _04738_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001110;
  assign _04739_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001101;
  assign _04740_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001100;
  assign _04741_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001011;
  assign _04742_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001010;
  assign _04743_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001001;
  assign _04744_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1001000;
  assign _04745_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000111;
  assign _04746_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000110;
  assign _04747_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000101;
  assign _04748_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000100;
  assign _04749_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000011;
  assign _04750_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000010;
  assign _04751_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000001;
  assign _04752_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 7'b1000000;
  assign _04753_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111111;
  assign _04754_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111110;
  assign _04755_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111101;
  assign _04756_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111100;
  assign _04757_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111011;
  assign _04758_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111010;
  assign _04759_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111001;
  assign _04760_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b111000;
  assign _04761_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110111;
  assign _04762_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110110;
  assign _04763_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110101;
  assign _04764_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110100;
  assign _04765_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110011;
  assign _04766_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110010;
  assign _04767_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110001;
  assign _04768_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b110000;
  assign _04769_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101111;
  assign _04770_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101110;
  assign _04771_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101101;
  assign _04772_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101100;
  assign _04773_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101011;
  assign _04774_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101010;
  assign _04775_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101001;
  assign _04776_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b101000;
  assign _04777_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100111;
  assign _04778_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100110;
  assign _04779_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100101;
  assign _04780_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100100;
  assign _04781_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100011;
  assign _04782_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100010;
  assign _04783_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100001;
  assign _04784_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 6'b100000;
  assign _04785_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11111;
  assign _04786_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11110;
  assign _04787_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11101;
  assign _04788_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11100;
  assign _04789_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11011;
  assign _04790_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11010;
  assign _04791_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11001;
  assign _04792_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b11000;
  assign _04793_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10111;
  assign _04794_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10110;
  assign _04795_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10101;
  assign _04796_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10100;
  assign _04797_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10011;
  assign _04798_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10010;
  assign _04799_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10001;
  assign _04800_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 5'b10000;
  assign _04801_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1111;
  assign _04802_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1110;
  assign _04803_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1101;
  assign _04804_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1100;
  assign _04805_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1011;
  assign _04806_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1010;
  assign _04807_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1001;
  assign _04808_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 4'b1000;
  assign _04809_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 3'b111;
  assign _04810_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 3'b110;
  assign _04811_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 3'b101;
  assign _04812_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 3'b100;
  assign _04813_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 2'b11;
  assign _04814_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 2'b10;
  assign _04815_ = vec_sum_091_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8805" *) 1'b1;
  function [7:0] _14243_;
    input [7:0] a;
    input [727:0] b;
    input [90:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *)
    (* parallel_case *)
    casez (s)
      91'b??????????????????????????????????????????????????????????????????????????????????????????1:
        _14243_ = b[7:0];
      91'b?????????????????????????????????????????????????????????????????????????????????????????1?:
        _14243_ = b[15:8];
      91'b????????????????????????????????????????????????????????????????????????????????????????1??:
        _14243_ = b[23:16];
      91'b???????????????????????????????????????????????????????????????????????????????????????1???:
        _14243_ = b[31:24];
      91'b??????????????????????????????????????????????????????????????????????????????????????1????:
        _14243_ = b[39:32];
      91'b?????????????????????????????????????????????????????????????????????????????????????1?????:
        _14243_ = b[47:40];
      91'b????????????????????????????????????????????????????????????????????????????????????1??????:
        _14243_ = b[55:48];
      91'b???????????????????????????????????????????????????????????????????????????????????1???????:
        _14243_ = b[63:56];
      91'b??????????????????????????????????????????????????????????????????????????????????1????????:
        _14243_ = b[71:64];
      91'b?????????????????????????????????????????????????????????????????????????????????1?????????:
        _14243_ = b[79:72];
      91'b????????????????????????????????????????????????????????????????????????????????1??????????:
        _14243_ = b[87:80];
      91'b???????????????????????????????????????????????????????????????????????????????1???????????:
        _14243_ = b[95:88];
      91'b??????????????????????????????????????????????????????????????????????????????1????????????:
        _14243_ = b[103:96];
      91'b?????????????????????????????????????????????????????????????????????????????1?????????????:
        _14243_ = b[111:104];
      91'b????????????????????????????????????????????????????????????????????????????1??????????????:
        _14243_ = b[119:112];
      91'b???????????????????????????????????????????????????????????????????????????1???????????????:
        _14243_ = b[127:120];
      91'b??????????????????????????????????????????????????????????????????????????1????????????????:
        _14243_ = b[135:128];
      91'b?????????????????????????????????????????????????????????????????????????1?????????????????:
        _14243_ = b[143:136];
      91'b????????????????????????????????????????????????????????????????????????1??????????????????:
        _14243_ = b[151:144];
      91'b???????????????????????????????????????????????????????????????????????1???????????????????:
        _14243_ = b[159:152];
      91'b??????????????????????????????????????????????????????????????????????1????????????????????:
        _14243_ = b[167:160];
      91'b?????????????????????????????????????????????????????????????????????1?????????????????????:
        _14243_ = b[175:168];
      91'b????????????????????????????????????????????????????????????????????1??????????????????????:
        _14243_ = b[183:176];
      91'b???????????????????????????????????????????????????????????????????1???????????????????????:
        _14243_ = b[191:184];
      91'b??????????????????????????????????????????????????????????????????1????????????????????????:
        _14243_ = b[199:192];
      91'b?????????????????????????????????????????????????????????????????1?????????????????????????:
        _14243_ = b[207:200];
      91'b????????????????????????????????????????????????????????????????1??????????????????????????:
        _14243_ = b[215:208];
      91'b???????????????????????????????????????????????????????????????1???????????????????????????:
        _14243_ = b[223:216];
      91'b??????????????????????????????????????????????????????????????1????????????????????????????:
        _14243_ = b[231:224];
      91'b?????????????????????????????????????????????????????????????1?????????????????????????????:
        _14243_ = b[239:232];
      91'b????????????????????????????????????????????????????????????1??????????????????????????????:
        _14243_ = b[247:240];
      91'b???????????????????????????????????????????????????????????1???????????????????????????????:
        _14243_ = b[255:248];
      91'b??????????????????????????????????????????????????????????1????????????????????????????????:
        _14243_ = b[263:256];
      91'b?????????????????????????????????????????????????????????1?????????????????????????????????:
        _14243_ = b[271:264];
      91'b????????????????????????????????????????????????????????1??????????????????????????????????:
        _14243_ = b[279:272];
      91'b???????????????????????????????????????????????????????1???????????????????????????????????:
        _14243_ = b[287:280];
      91'b??????????????????????????????????????????????????????1????????????????????????????????????:
        _14243_ = b[295:288];
      91'b?????????????????????????????????????????????????????1?????????????????????????????????????:
        _14243_ = b[303:296];
      91'b????????????????????????????????????????????????????1??????????????????????????????????????:
        _14243_ = b[311:304];
      91'b???????????????????????????????????????????????????1???????????????????????????????????????:
        _14243_ = b[319:312];
      91'b??????????????????????????????????????????????????1????????????????????????????????????????:
        _14243_ = b[327:320];
      91'b?????????????????????????????????????????????????1?????????????????????????????????????????:
        _14243_ = b[335:328];
      91'b????????????????????????????????????????????????1??????????????????????????????????????????:
        _14243_ = b[343:336];
      91'b???????????????????????????????????????????????1???????????????????????????????????????????:
        _14243_ = b[351:344];
      91'b??????????????????????????????????????????????1????????????????????????????????????????????:
        _14243_ = b[359:352];
      91'b?????????????????????????????????????????????1?????????????????????????????????????????????:
        _14243_ = b[367:360];
      91'b????????????????????????????????????????????1??????????????????????????????????????????????:
        _14243_ = b[375:368];
      91'b???????????????????????????????????????????1???????????????????????????????????????????????:
        _14243_ = b[383:376];
      91'b??????????????????????????????????????????1????????????????????????????????????????????????:
        _14243_ = b[391:384];
      91'b?????????????????????????????????????????1?????????????????????????????????????????????????:
        _14243_ = b[399:392];
      91'b????????????????????????????????????????1??????????????????????????????????????????????????:
        _14243_ = b[407:400];
      91'b???????????????????????????????????????1???????????????????????????????????????????????????:
        _14243_ = b[415:408];
      91'b??????????????????????????????????????1????????????????????????????????????????????????????:
        _14243_ = b[423:416];
      91'b?????????????????????????????????????1?????????????????????????????????????????????????????:
        _14243_ = b[431:424];
      91'b????????????????????????????????????1??????????????????????????????????????????????????????:
        _14243_ = b[439:432];
      91'b???????????????????????????????????1???????????????????????????????????????????????????????:
        _14243_ = b[447:440];
      91'b??????????????????????????????????1????????????????????????????????????????????????????????:
        _14243_ = b[455:448];
      91'b?????????????????????????????????1?????????????????????????????????????????????????????????:
        _14243_ = b[463:456];
      91'b????????????????????????????????1??????????????????????????????????????????????????????????:
        _14243_ = b[471:464];
      91'b???????????????????????????????1???????????????????????????????????????????????????????????:
        _14243_ = b[479:472];
      91'b??????????????????????????????1????????????????????????????????????????????????????????????:
        _14243_ = b[487:480];
      91'b?????????????????????????????1?????????????????????????????????????????????????????????????:
        _14243_ = b[495:488];
      91'b????????????????????????????1??????????????????????????????????????????????????????????????:
        _14243_ = b[503:496];
      91'b???????????????????????????1???????????????????????????????????????????????????????????????:
        _14243_ = b[511:504];
      91'b??????????????????????????1????????????????????????????????????????????????????????????????:
        _14243_ = b[519:512];
      91'b?????????????????????????1?????????????????????????????????????????????????????????????????:
        _14243_ = b[527:520];
      91'b????????????????????????1??????????????????????????????????????????????????????????????????:
        _14243_ = b[535:528];
      91'b???????????????????????1???????????????????????????????????????????????????????????????????:
        _14243_ = b[543:536];
      91'b??????????????????????1????????????????????????????????????????????????????????????????????:
        _14243_ = b[551:544];
      91'b?????????????????????1?????????????????????????????????????????????????????????????????????:
        _14243_ = b[559:552];
      91'b????????????????????1??????????????????????????????????????????????????????????????????????:
        _14243_ = b[567:560];
      91'b???????????????????1???????????????????????????????????????????????????????????????????????:
        _14243_ = b[575:568];
      91'b??????????????????1????????????????????????????????????????????????????????????????????????:
        _14243_ = b[583:576];
      91'b?????????????????1?????????????????????????????????????????????????????????????????????????:
        _14243_ = b[591:584];
      91'b????????????????1??????????????????????????????????????????????????????????????????????????:
        _14243_ = b[599:592];
      91'b???????????????1???????????????????????????????????????????????????????????????????????????:
        _14243_ = b[607:600];
      91'b??????????????1????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[615:608];
      91'b?????????????1?????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[623:616];
      91'b????????????1??????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[631:624];
      91'b???????????1???????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[639:632];
      91'b??????????1????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[647:640];
      91'b?????????1?????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[655:648];
      91'b????????1??????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[663:656];
      91'b???????1???????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[671:664];
      91'b??????1????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[679:672];
      91'b?????1?????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[687:680];
      91'b????1??????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[695:688];
      91'b???1???????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[703:696];
      91'b??1????????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[711:704];
      91'b?1?????????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[719:712];
      91'b1??????????????????????????????????????????????????????????????????????????????????????????:
        _14243_ = b[727:720];
      default:
        _14243_ = a;
    endcase
  endfunction
  assign vec_data_090 = _14243_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712], data_d1[727:720] }, { _04906_, _04905_, _04904_, _04903_, _04902_, _04901_, _04900_, _04899_, _04898_, _04897_, _04896_, _04895_, _04894_, _04893_, _04892_, _04891_, _04890_, _04889_, _04888_, _04887_, _04886_, _04885_, _04884_, _04883_, _04882_, _04881_, _04880_, _04879_, _04878_, _04877_, _04876_, _04875_, _04874_, _04873_, _04872_, _04871_, _04870_, _04869_, _04868_, _04867_, _04866_, _04865_, _04864_, _04863_, _04862_, _04861_, _04860_, _04859_, _04858_, _04857_, _04856_, _04855_, _04854_, _04853_, _04852_, _04851_, _04850_, _04849_, _04848_, _04847_, _04846_, _04845_, _04844_, _04843_, _04842_, _04841_, _04840_, _04839_, _04838_, _04837_, _04836_, _04835_, _04834_, _04833_, _04832_, _04831_, _04830_, _04829_, _04828_, _04827_, _04826_, _04825_, _04824_, _04823_, _04822_, _04821_, _04820_, _04819_, _04818_, _04817_, _04816_ });
  assign _04816_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1011011;
  assign _04817_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1011010;
  assign _04818_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1011001;
  assign _04819_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1011000;
  assign _04820_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010111;
  assign _04821_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010110;
  assign _04822_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010101;
  assign _04823_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010100;
  assign _04824_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010011;
  assign _04825_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010010;
  assign _04826_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010001;
  assign _04827_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1010000;
  assign _04828_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001111;
  assign _04829_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001110;
  assign _04830_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001101;
  assign _04831_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001100;
  assign _04832_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001011;
  assign _04833_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001010;
  assign _04834_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001001;
  assign _04835_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1001000;
  assign _04836_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000111;
  assign _04837_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000110;
  assign _04838_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000101;
  assign _04839_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000100;
  assign _04840_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000011;
  assign _04841_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000010;
  assign _04842_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000001;
  assign _04843_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 7'b1000000;
  assign _04844_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111111;
  assign _04845_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111110;
  assign _04846_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111101;
  assign _04847_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111100;
  assign _04848_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111011;
  assign _04849_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111010;
  assign _04850_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111001;
  assign _04851_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b111000;
  assign _04852_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110111;
  assign _04853_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110110;
  assign _04854_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110101;
  assign _04855_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110100;
  assign _04856_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110011;
  assign _04857_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110010;
  assign _04858_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110001;
  assign _04859_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b110000;
  assign _04860_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101111;
  assign _04861_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101110;
  assign _04862_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101101;
  assign _04863_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101100;
  assign _04864_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101011;
  assign _04865_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101010;
  assign _04866_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101001;
  assign _04867_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b101000;
  assign _04868_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100111;
  assign _04869_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100110;
  assign _04870_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100101;
  assign _04871_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100100;
  assign _04872_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100011;
  assign _04873_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100010;
  assign _04874_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100001;
  assign _04875_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 6'b100000;
  assign _04876_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11111;
  assign _04877_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11110;
  assign _04878_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11101;
  assign _04879_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11100;
  assign _04880_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11011;
  assign _04881_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11010;
  assign _04882_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11001;
  assign _04883_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b11000;
  assign _04884_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10111;
  assign _04885_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10110;
  assign _04886_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10101;
  assign _04887_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10100;
  assign _04888_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10011;
  assign _04889_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10010;
  assign _04890_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10001;
  assign _04891_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 5'b10000;
  assign _04892_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1111;
  assign _04893_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1110;
  assign _04894_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1101;
  assign _04895_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1100;
  assign _04896_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1011;
  assign _04897_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1010;
  assign _04898_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1001;
  assign _04899_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 4'b1000;
  assign _04900_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 3'b111;
  assign _04901_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 3'b110;
  assign _04902_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 3'b101;
  assign _04903_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 3'b100;
  assign _04904_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 2'b11;
  assign _04905_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 2'b10;
  assign _04906_ = vec_sum_090_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8706" *) 1'b1;
  function [7:0] _14335_;
    input [7:0] a;
    input [719:0] b;
    input [89:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *)
    (* parallel_case *)
    casez (s)
      90'b?????????????????????????????????????????????????????????????????????????????????????????1:
        _14335_ = b[7:0];
      90'b????????????????????????????????????????????????????????????????????????????????????????1?:
        _14335_ = b[15:8];
      90'b???????????????????????????????????????????????????????????????????????????????????????1??:
        _14335_ = b[23:16];
      90'b??????????????????????????????????????????????????????????????????????????????????????1???:
        _14335_ = b[31:24];
      90'b?????????????????????????????????????????????????????????????????????????????????????1????:
        _14335_ = b[39:32];
      90'b????????????????????????????????????????????????????????????????????????????????????1?????:
        _14335_ = b[47:40];
      90'b???????????????????????????????????????????????????????????????????????????????????1??????:
        _14335_ = b[55:48];
      90'b??????????????????????????????????????????????????????????????????????????????????1???????:
        _14335_ = b[63:56];
      90'b?????????????????????????????????????????????????????????????????????????????????1????????:
        _14335_ = b[71:64];
      90'b????????????????????????????????????????????????????????????????????????????????1?????????:
        _14335_ = b[79:72];
      90'b???????????????????????????????????????????????????????????????????????????????1??????????:
        _14335_ = b[87:80];
      90'b??????????????????????????????????????????????????????????????????????????????1???????????:
        _14335_ = b[95:88];
      90'b?????????????????????????????????????????????????????????????????????????????1????????????:
        _14335_ = b[103:96];
      90'b????????????????????????????????????????????????????????????????????????????1?????????????:
        _14335_ = b[111:104];
      90'b???????????????????????????????????????????????????????????????????????????1??????????????:
        _14335_ = b[119:112];
      90'b??????????????????????????????????????????????????????????????????????????1???????????????:
        _14335_ = b[127:120];
      90'b?????????????????????????????????????????????????????????????????????????1????????????????:
        _14335_ = b[135:128];
      90'b????????????????????????????????????????????????????????????????????????1?????????????????:
        _14335_ = b[143:136];
      90'b???????????????????????????????????????????????????????????????????????1??????????????????:
        _14335_ = b[151:144];
      90'b??????????????????????????????????????????????????????????????????????1???????????????????:
        _14335_ = b[159:152];
      90'b?????????????????????????????????????????????????????????????????????1????????????????????:
        _14335_ = b[167:160];
      90'b????????????????????????????????????????????????????????????????????1?????????????????????:
        _14335_ = b[175:168];
      90'b???????????????????????????????????????????????????????????????????1??????????????????????:
        _14335_ = b[183:176];
      90'b??????????????????????????????????????????????????????????????????1???????????????????????:
        _14335_ = b[191:184];
      90'b?????????????????????????????????????????????????????????????????1????????????????????????:
        _14335_ = b[199:192];
      90'b????????????????????????????????????????????????????????????????1?????????????????????????:
        _14335_ = b[207:200];
      90'b???????????????????????????????????????????????????????????????1??????????????????????????:
        _14335_ = b[215:208];
      90'b??????????????????????????????????????????????????????????????1???????????????????????????:
        _14335_ = b[223:216];
      90'b?????????????????????????????????????????????????????????????1????????????????????????????:
        _14335_ = b[231:224];
      90'b????????????????????????????????????????????????????????????1?????????????????????????????:
        _14335_ = b[239:232];
      90'b???????????????????????????????????????????????????????????1??????????????????????????????:
        _14335_ = b[247:240];
      90'b??????????????????????????????????????????????????????????1???????????????????????????????:
        _14335_ = b[255:248];
      90'b?????????????????????????????????????????????????????????1????????????????????????????????:
        _14335_ = b[263:256];
      90'b????????????????????????????????????????????????????????1?????????????????????????????????:
        _14335_ = b[271:264];
      90'b???????????????????????????????????????????????????????1??????????????????????????????????:
        _14335_ = b[279:272];
      90'b??????????????????????????????????????????????????????1???????????????????????????????????:
        _14335_ = b[287:280];
      90'b?????????????????????????????????????????????????????1????????????????????????????????????:
        _14335_ = b[295:288];
      90'b????????????????????????????????????????????????????1?????????????????????????????????????:
        _14335_ = b[303:296];
      90'b???????????????????????????????????????????????????1??????????????????????????????????????:
        _14335_ = b[311:304];
      90'b??????????????????????????????????????????????????1???????????????????????????????????????:
        _14335_ = b[319:312];
      90'b?????????????????????????????????????????????????1????????????????????????????????????????:
        _14335_ = b[327:320];
      90'b????????????????????????????????????????????????1?????????????????????????????????????????:
        _14335_ = b[335:328];
      90'b???????????????????????????????????????????????1??????????????????????????????????????????:
        _14335_ = b[343:336];
      90'b??????????????????????????????????????????????1???????????????????????????????????????????:
        _14335_ = b[351:344];
      90'b?????????????????????????????????????????????1????????????????????????????????????????????:
        _14335_ = b[359:352];
      90'b????????????????????????????????????????????1?????????????????????????????????????????????:
        _14335_ = b[367:360];
      90'b???????????????????????????????????????????1??????????????????????????????????????????????:
        _14335_ = b[375:368];
      90'b??????????????????????????????????????????1???????????????????????????????????????????????:
        _14335_ = b[383:376];
      90'b?????????????????????????????????????????1????????????????????????????????????????????????:
        _14335_ = b[391:384];
      90'b????????????????????????????????????????1?????????????????????????????????????????????????:
        _14335_ = b[399:392];
      90'b???????????????????????????????????????1??????????????????????????????????????????????????:
        _14335_ = b[407:400];
      90'b??????????????????????????????????????1???????????????????????????????????????????????????:
        _14335_ = b[415:408];
      90'b?????????????????????????????????????1????????????????????????????????????????????????????:
        _14335_ = b[423:416];
      90'b????????????????????????????????????1?????????????????????????????????????????????????????:
        _14335_ = b[431:424];
      90'b???????????????????????????????????1??????????????????????????????????????????????????????:
        _14335_ = b[439:432];
      90'b??????????????????????????????????1???????????????????????????????????????????????????????:
        _14335_ = b[447:440];
      90'b?????????????????????????????????1????????????????????????????????????????????????????????:
        _14335_ = b[455:448];
      90'b????????????????????????????????1?????????????????????????????????????????????????????????:
        _14335_ = b[463:456];
      90'b???????????????????????????????1??????????????????????????????????????????????????????????:
        _14335_ = b[471:464];
      90'b??????????????????????????????1???????????????????????????????????????????????????????????:
        _14335_ = b[479:472];
      90'b?????????????????????????????1????????????????????????????????????????????????????????????:
        _14335_ = b[487:480];
      90'b????????????????????????????1?????????????????????????????????????????????????????????????:
        _14335_ = b[495:488];
      90'b???????????????????????????1??????????????????????????????????????????????????????????????:
        _14335_ = b[503:496];
      90'b??????????????????????????1???????????????????????????????????????????????????????????????:
        _14335_ = b[511:504];
      90'b?????????????????????????1????????????????????????????????????????????????????????????????:
        _14335_ = b[519:512];
      90'b????????????????????????1?????????????????????????????????????????????????????????????????:
        _14335_ = b[527:520];
      90'b???????????????????????1??????????????????????????????????????????????????????????????????:
        _14335_ = b[535:528];
      90'b??????????????????????1???????????????????????????????????????????????????????????????????:
        _14335_ = b[543:536];
      90'b?????????????????????1????????????????????????????????????????????????????????????????????:
        _14335_ = b[551:544];
      90'b????????????????????1?????????????????????????????????????????????????????????????????????:
        _14335_ = b[559:552];
      90'b???????????????????1??????????????????????????????????????????????????????????????????????:
        _14335_ = b[567:560];
      90'b??????????????????1???????????????????????????????????????????????????????????????????????:
        _14335_ = b[575:568];
      90'b?????????????????1????????????????????????????????????????????????????????????????????????:
        _14335_ = b[583:576];
      90'b????????????????1?????????????????????????????????????????????????????????????????????????:
        _14335_ = b[591:584];
      90'b???????????????1??????????????????????????????????????????????????????????????????????????:
        _14335_ = b[599:592];
      90'b??????????????1???????????????????????????????????????????????????????????????????????????:
        _14335_ = b[607:600];
      90'b?????????????1????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[615:608];
      90'b????????????1?????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[623:616];
      90'b???????????1??????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[631:624];
      90'b??????????1???????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[639:632];
      90'b?????????1????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[647:640];
      90'b????????1?????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[655:648];
      90'b???????1??????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[663:656];
      90'b??????1???????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[671:664];
      90'b?????1????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[679:672];
      90'b????1?????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[687:680];
      90'b???1??????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[695:688];
      90'b??1???????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[703:696];
      90'b?1????????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[711:704];
      90'b1?????????????????????????????????????????????????????????????????????????????????????????:
        _14335_ = b[719:712];
      default:
        _14335_ = a;
    endcase
  endfunction
  assign vec_data_089 = _14335_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704], data_d1[719:712] }, { _04996_, _04995_, _04994_, _04993_, _04992_, _04991_, _04990_, _04989_, _04988_, _04987_, _04986_, _04985_, _04984_, _04983_, _04982_, _04981_, _04980_, _04979_, _04978_, _04977_, _04976_, _04975_, _04974_, _04973_, _04972_, _04971_, _04970_, _04969_, _04968_, _04967_, _04966_, _04965_, _04964_, _04963_, _04962_, _04961_, _04960_, _04959_, _04958_, _04957_, _04956_, _04955_, _04954_, _04953_, _04952_, _04951_, _04950_, _04949_, _04948_, _04947_, _04946_, _04945_, _04944_, _04943_, _04942_, _04941_, _04940_, _04939_, _04938_, _04937_, _04936_, _04935_, _04934_, _04933_, _04932_, _04931_, _04930_, _04929_, _04928_, _04927_, _04926_, _04925_, _04924_, _04923_, _04922_, _04921_, _04920_, _04919_, _04918_, _04917_, _04916_, _04915_, _04914_, _04913_, _04912_, _04911_, _04910_, _04909_, _04908_, _04907_ });
  assign _04907_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1011010;
  assign _04908_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1011001;
  assign _04909_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1011000;
  assign _04910_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010111;
  assign _04911_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010110;
  assign _04912_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010101;
  assign _04913_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010100;
  assign _04914_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010011;
  assign _04915_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010010;
  assign _04916_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010001;
  assign _04917_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1010000;
  assign _04918_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001111;
  assign _04919_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001110;
  assign _04920_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001101;
  assign _04921_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001100;
  assign _04922_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001011;
  assign _04923_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001010;
  assign _04924_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001001;
  assign _04925_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1001000;
  assign _04926_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000111;
  assign _04927_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000110;
  assign _04928_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000101;
  assign _04929_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000100;
  assign _04930_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000011;
  assign _04931_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000010;
  assign _04932_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000001;
  assign _04933_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 7'b1000000;
  assign _04934_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111111;
  assign _04935_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111110;
  assign _04936_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111101;
  assign _04937_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111100;
  assign _04938_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111011;
  assign _04939_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111010;
  assign _04940_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111001;
  assign _04941_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b111000;
  assign _04942_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110111;
  assign _04943_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110110;
  assign _04944_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110101;
  assign _04945_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110100;
  assign _04946_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110011;
  assign _04947_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110010;
  assign _04948_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110001;
  assign _04949_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b110000;
  assign _04950_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101111;
  assign _04951_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101110;
  assign _04952_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101101;
  assign _04953_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101100;
  assign _04954_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101011;
  assign _04955_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101010;
  assign _04956_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101001;
  assign _04957_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b101000;
  assign _04958_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100111;
  assign _04959_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100110;
  assign _04960_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100101;
  assign _04961_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100100;
  assign _04962_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100011;
  assign _04963_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100010;
  assign _04964_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100001;
  assign _04965_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 6'b100000;
  assign _04966_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11111;
  assign _04967_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11110;
  assign _04968_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11101;
  assign _04969_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11100;
  assign _04970_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11011;
  assign _04971_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11010;
  assign _04972_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11001;
  assign _04973_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b11000;
  assign _04974_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10111;
  assign _04975_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8630|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10110;
  assign _04976_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8629|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10101;
  assign _04977_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8628|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10100;
  assign _04978_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10011;
  assign _04979_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10010;
  assign _04980_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10001;
  assign _04981_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 5'b10000;
  assign _04982_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1111;
  assign _04983_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1110;
  assign _04984_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1101;
  assign _04985_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1100;
  assign _04986_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1011;
  assign _04987_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1010;
  assign _04988_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1001;
  assign _04989_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 4'b1000;
  assign _04990_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 3'b111;
  assign _04991_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 3'b110;
  assign _04992_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 3'b101;
  assign _04993_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 3'b100;
  assign _04994_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 2'b11;
  assign _04995_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 2'b10;
  assign _04996_ = vec_sum_089_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8608" *) 1'b1;
  function [7:0] _14426_;
    input [7:0] a;
    input [711:0] b;
    input [88:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *)
    (* parallel_case *)
    casez (s)
      89'b????????????????????????????????????????????????????????????????????????????????????????1:
        _14426_ = b[7:0];
      89'b???????????????????????????????????????????????????????????????????????????????????????1?:
        _14426_ = b[15:8];
      89'b??????????????????????????????????????????????????????????????????????????????????????1??:
        _14426_ = b[23:16];
      89'b?????????????????????????????????????????????????????????????????????????????????????1???:
        _14426_ = b[31:24];
      89'b????????????????????????????????????????????????????????????????????????????????????1????:
        _14426_ = b[39:32];
      89'b???????????????????????????????????????????????????????????????????????????????????1?????:
        _14426_ = b[47:40];
      89'b??????????????????????????????????????????????????????????????????????????????????1??????:
        _14426_ = b[55:48];
      89'b?????????????????????????????????????????????????????????????????????????????????1???????:
        _14426_ = b[63:56];
      89'b????????????????????????????????????????????????????????????????????????????????1????????:
        _14426_ = b[71:64];
      89'b???????????????????????????????????????????????????????????????????????????????1?????????:
        _14426_ = b[79:72];
      89'b??????????????????????????????????????????????????????????????????????????????1??????????:
        _14426_ = b[87:80];
      89'b?????????????????????????????????????????????????????????????????????????????1???????????:
        _14426_ = b[95:88];
      89'b????????????????????????????????????????????????????????????????????????????1????????????:
        _14426_ = b[103:96];
      89'b???????????????????????????????????????????????????????????????????????????1?????????????:
        _14426_ = b[111:104];
      89'b??????????????????????????????????????????????????????????????????????????1??????????????:
        _14426_ = b[119:112];
      89'b?????????????????????????????????????????????????????????????????????????1???????????????:
        _14426_ = b[127:120];
      89'b????????????????????????????????????????????????????????????????????????1????????????????:
        _14426_ = b[135:128];
      89'b???????????????????????????????????????????????????????????????????????1?????????????????:
        _14426_ = b[143:136];
      89'b??????????????????????????????????????????????????????????????????????1??????????????????:
        _14426_ = b[151:144];
      89'b?????????????????????????????????????????????????????????????????????1???????????????????:
        _14426_ = b[159:152];
      89'b????????????????????????????????????????????????????????????????????1????????????????????:
        _14426_ = b[167:160];
      89'b???????????????????????????????????????????????????????????????????1?????????????????????:
        _14426_ = b[175:168];
      89'b??????????????????????????????????????????????????????????????????1??????????????????????:
        _14426_ = b[183:176];
      89'b?????????????????????????????????????????????????????????????????1???????????????????????:
        _14426_ = b[191:184];
      89'b????????????????????????????????????????????????????????????????1????????????????????????:
        _14426_ = b[199:192];
      89'b???????????????????????????????????????????????????????????????1?????????????????????????:
        _14426_ = b[207:200];
      89'b??????????????????????????????????????????????????????????????1??????????????????????????:
        _14426_ = b[215:208];
      89'b?????????????????????????????????????????????????????????????1???????????????????????????:
        _14426_ = b[223:216];
      89'b????????????????????????????????????????????????????????????1????????????????????????????:
        _14426_ = b[231:224];
      89'b???????????????????????????????????????????????????????????1?????????????????????????????:
        _14426_ = b[239:232];
      89'b??????????????????????????????????????????????????????????1??????????????????????????????:
        _14426_ = b[247:240];
      89'b?????????????????????????????????????????????????????????1???????????????????????????????:
        _14426_ = b[255:248];
      89'b????????????????????????????????????????????????????????1????????????????????????????????:
        _14426_ = b[263:256];
      89'b???????????????????????????????????????????????????????1?????????????????????????????????:
        _14426_ = b[271:264];
      89'b??????????????????????????????????????????????????????1??????????????????????????????????:
        _14426_ = b[279:272];
      89'b?????????????????????????????????????????????????????1???????????????????????????????????:
        _14426_ = b[287:280];
      89'b????????????????????????????????????????????????????1????????????????????????????????????:
        _14426_ = b[295:288];
      89'b???????????????????????????????????????????????????1?????????????????????????????????????:
        _14426_ = b[303:296];
      89'b??????????????????????????????????????????????????1??????????????????????????????????????:
        _14426_ = b[311:304];
      89'b?????????????????????????????????????????????????1???????????????????????????????????????:
        _14426_ = b[319:312];
      89'b????????????????????????????????????????????????1????????????????????????????????????????:
        _14426_ = b[327:320];
      89'b???????????????????????????????????????????????1?????????????????????????????????????????:
        _14426_ = b[335:328];
      89'b??????????????????????????????????????????????1??????????????????????????????????????????:
        _14426_ = b[343:336];
      89'b?????????????????????????????????????????????1???????????????????????????????????????????:
        _14426_ = b[351:344];
      89'b????????????????????????????????????????????1????????????????????????????????????????????:
        _14426_ = b[359:352];
      89'b???????????????????????????????????????????1?????????????????????????????????????????????:
        _14426_ = b[367:360];
      89'b??????????????????????????????????????????1??????????????????????????????????????????????:
        _14426_ = b[375:368];
      89'b?????????????????????????????????????????1???????????????????????????????????????????????:
        _14426_ = b[383:376];
      89'b????????????????????????????????????????1????????????????????????????????????????????????:
        _14426_ = b[391:384];
      89'b???????????????????????????????????????1?????????????????????????????????????????????????:
        _14426_ = b[399:392];
      89'b??????????????????????????????????????1??????????????????????????????????????????????????:
        _14426_ = b[407:400];
      89'b?????????????????????????????????????1???????????????????????????????????????????????????:
        _14426_ = b[415:408];
      89'b????????????????????????????????????1????????????????????????????????????????????????????:
        _14426_ = b[423:416];
      89'b???????????????????????????????????1?????????????????????????????????????????????????????:
        _14426_ = b[431:424];
      89'b??????????????????????????????????1??????????????????????????????????????????????????????:
        _14426_ = b[439:432];
      89'b?????????????????????????????????1???????????????????????????????????????????????????????:
        _14426_ = b[447:440];
      89'b????????????????????????????????1????????????????????????????????????????????????????????:
        _14426_ = b[455:448];
      89'b???????????????????????????????1?????????????????????????????????????????????????????????:
        _14426_ = b[463:456];
      89'b??????????????????????????????1??????????????????????????????????????????????????????????:
        _14426_ = b[471:464];
      89'b?????????????????????????????1???????????????????????????????????????????????????????????:
        _14426_ = b[479:472];
      89'b????????????????????????????1????????????????????????????????????????????????????????????:
        _14426_ = b[487:480];
      89'b???????????????????????????1?????????????????????????????????????????????????????????????:
        _14426_ = b[495:488];
      89'b??????????????????????????1??????????????????????????????????????????????????????????????:
        _14426_ = b[503:496];
      89'b?????????????????????????1???????????????????????????????????????????????????????????????:
        _14426_ = b[511:504];
      89'b????????????????????????1????????????????????????????????????????????????????????????????:
        _14426_ = b[519:512];
      89'b???????????????????????1?????????????????????????????????????????????????????????????????:
        _14426_ = b[527:520];
      89'b??????????????????????1??????????????????????????????????????????????????????????????????:
        _14426_ = b[535:528];
      89'b?????????????????????1???????????????????????????????????????????????????????????????????:
        _14426_ = b[543:536];
      89'b????????????????????1????????????????????????????????????????????????????????????????????:
        _14426_ = b[551:544];
      89'b???????????????????1?????????????????????????????????????????????????????????????????????:
        _14426_ = b[559:552];
      89'b??????????????????1??????????????????????????????????????????????????????????????????????:
        _14426_ = b[567:560];
      89'b?????????????????1???????????????????????????????????????????????????????????????????????:
        _14426_ = b[575:568];
      89'b????????????????1????????????????????????????????????????????????????????????????????????:
        _14426_ = b[583:576];
      89'b???????????????1?????????????????????????????????????????????????????????????????????????:
        _14426_ = b[591:584];
      89'b??????????????1??????????????????????????????????????????????????????????????????????????:
        _14426_ = b[599:592];
      89'b?????????????1???????????????????????????????????????????????????????????????????????????:
        _14426_ = b[607:600];
      89'b????????????1????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[615:608];
      89'b???????????1?????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[623:616];
      89'b??????????1??????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[631:624];
      89'b?????????1???????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[639:632];
      89'b????????1????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[647:640];
      89'b???????1?????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[655:648];
      89'b??????1??????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[663:656];
      89'b?????1???????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[671:664];
      89'b????1????????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[679:672];
      89'b???1?????????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[687:680];
      89'b??1??????????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[695:688];
      89'b?1???????????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[703:696];
      89'b1????????????????????????????????????????????????????????????????????????????????????????:
        _14426_ = b[711:704];
      default:
        _14426_ = a;
    endcase
  endfunction
  assign vec_data_088 = _14426_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696], data_d1[711:704] }, { _05085_, _05084_, _05083_, _05082_, _05081_, _05080_, _05079_, _05078_, _05077_, _05076_, _05075_, _05074_, _05073_, _05072_, _05071_, _05070_, _05069_, _05068_, _05067_, _05066_, _05065_, _05064_, _05063_, _05062_, _05061_, _05060_, _05059_, _05058_, _05057_, _05056_, _05055_, _05054_, _05053_, _05052_, _05051_, _05050_, _05049_, _05048_, _05047_, _05046_, _05045_, _05044_, _05043_, _05042_, _05041_, _05040_, _05039_, _05038_, _05037_, _05036_, _05035_, _05034_, _05033_, _05032_, _05031_, _05030_, _05029_, _05028_, _05027_, _05026_, _05025_, _05024_, _05023_, _05022_, _05021_, _05020_, _05019_, _05018_, _05017_, _05016_, _05015_, _05014_, _05013_, _05012_, _05011_, _05010_, _05009_, _05008_, _05007_, _05006_, _05005_, _05004_, _05003_, _05002_, _05001_, _05000_, _04999_, _04998_, _04997_ });
  assign _04997_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1011001;
  assign _04998_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1011000;
  assign _04999_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010111;
  assign _05000_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010110;
  assign _05001_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010101;
  assign _05002_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010100;
  assign _05003_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010011;
  assign _05004_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010010;
  assign _05005_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010001;
  assign _05006_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1010000;
  assign _05007_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001111;
  assign _05008_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001110;
  assign _05009_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001101;
  assign _05010_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001100;
  assign _05011_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001011;
  assign _05012_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001010;
  assign _05013_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001001;
  assign _05014_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1001000;
  assign _05015_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000111;
  assign _05016_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000110;
  assign _05017_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000101;
  assign _05018_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000100;
  assign _05019_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000011;
  assign _05020_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000010;
  assign _05021_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000001;
  assign _05022_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 7'b1000000;
  assign _05023_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111111;
  assign _05024_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111110;
  assign _05025_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111101;
  assign _05026_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111100;
  assign _05027_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111011;
  assign _05028_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111010;
  assign _05029_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111001;
  assign _05030_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b111000;
  assign _05031_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110111;
  assign _05032_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110110;
  assign _05033_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110101;
  assign _05034_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110100;
  assign _05035_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110011;
  assign _05036_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110010;
  assign _05037_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110001;
  assign _05038_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b110000;
  assign _05039_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101111;
  assign _05040_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101110;
  assign _05041_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101101;
  assign _05042_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101100;
  assign _05043_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101011;
  assign _05044_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101010;
  assign _05045_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101001;
  assign _05046_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b101000;
  assign _05047_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100111;
  assign _05048_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100110;
  assign _05049_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100101;
  assign _05050_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100100;
  assign _05051_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100011;
  assign _05052_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100010;
  assign _05053_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100001;
  assign _05054_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 6'b100000;
  assign _05055_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11111;
  assign _05056_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11110;
  assign _05057_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11101;
  assign _05058_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11100;
  assign _05059_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11011;
  assign _05060_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11010;
  assign _05061_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11001;
  assign _05062_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b11000;
  assign _05063_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10111;
  assign _05064_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10110;
  assign _05065_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10101;
  assign _05066_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10100;
  assign _05067_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10011;
  assign _05068_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10010;
  assign _05069_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10001;
  assign _05070_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 5'b10000;
  assign _05071_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1111;
  assign _05072_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1110;
  assign _05073_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1101;
  assign _05074_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1100;
  assign _05075_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1011;
  assign _05076_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1010;
  assign _05077_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1001;
  assign _05078_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 4'b1000;
  assign _05079_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 3'b111;
  assign _05080_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 3'b110;
  assign _05081_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 3'b101;
  assign _05082_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 3'b100;
  assign _05083_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 2'b11;
  assign _05084_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 2'b10;
  assign _05085_ = vec_sum_088_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8511" *) 1'b1;
  function [7:0] _14516_;
    input [7:0] a;
    input [703:0] b;
    input [87:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *)
    (* parallel_case *)
    casez (s)
      88'b???????????????????????????????????????????????????????????????????????????????????????1:
        _14516_ = b[7:0];
      88'b??????????????????????????????????????????????????????????????????????????????????????1?:
        _14516_ = b[15:8];
      88'b?????????????????????????????????????????????????????????????????????????????????????1??:
        _14516_ = b[23:16];
      88'b????????????????????????????????????????????????????????????????????????????????????1???:
        _14516_ = b[31:24];
      88'b???????????????????????????????????????????????????????????????????????????????????1????:
        _14516_ = b[39:32];
      88'b??????????????????????????????????????????????????????????????????????????????????1?????:
        _14516_ = b[47:40];
      88'b?????????????????????????????????????????????????????????????????????????????????1??????:
        _14516_ = b[55:48];
      88'b????????????????????????????????????????????????????????????????????????????????1???????:
        _14516_ = b[63:56];
      88'b???????????????????????????????????????????????????????????????????????????????1????????:
        _14516_ = b[71:64];
      88'b??????????????????????????????????????????????????????????????????????????????1?????????:
        _14516_ = b[79:72];
      88'b?????????????????????????????????????????????????????????????????????????????1??????????:
        _14516_ = b[87:80];
      88'b????????????????????????????????????????????????????????????????????????????1???????????:
        _14516_ = b[95:88];
      88'b???????????????????????????????????????????????????????????????????????????1????????????:
        _14516_ = b[103:96];
      88'b??????????????????????????????????????????????????????????????????????????1?????????????:
        _14516_ = b[111:104];
      88'b?????????????????????????????????????????????????????????????????????????1??????????????:
        _14516_ = b[119:112];
      88'b????????????????????????????????????????????????????????????????????????1???????????????:
        _14516_ = b[127:120];
      88'b???????????????????????????????????????????????????????????????????????1????????????????:
        _14516_ = b[135:128];
      88'b??????????????????????????????????????????????????????????????????????1?????????????????:
        _14516_ = b[143:136];
      88'b?????????????????????????????????????????????????????????????????????1??????????????????:
        _14516_ = b[151:144];
      88'b????????????????????????????????????????????????????????????????????1???????????????????:
        _14516_ = b[159:152];
      88'b???????????????????????????????????????????????????????????????????1????????????????????:
        _14516_ = b[167:160];
      88'b??????????????????????????????????????????????????????????????????1?????????????????????:
        _14516_ = b[175:168];
      88'b?????????????????????????????????????????????????????????????????1??????????????????????:
        _14516_ = b[183:176];
      88'b????????????????????????????????????????????????????????????????1???????????????????????:
        _14516_ = b[191:184];
      88'b???????????????????????????????????????????????????????????????1????????????????????????:
        _14516_ = b[199:192];
      88'b??????????????????????????????????????????????????????????????1?????????????????????????:
        _14516_ = b[207:200];
      88'b?????????????????????????????????????????????????????????????1??????????????????????????:
        _14516_ = b[215:208];
      88'b????????????????????????????????????????????????????????????1???????????????????????????:
        _14516_ = b[223:216];
      88'b???????????????????????????????????????????????????????????1????????????????????????????:
        _14516_ = b[231:224];
      88'b??????????????????????????????????????????????????????????1?????????????????????????????:
        _14516_ = b[239:232];
      88'b?????????????????????????????????????????????????????????1??????????????????????????????:
        _14516_ = b[247:240];
      88'b????????????????????????????????????????????????????????1???????????????????????????????:
        _14516_ = b[255:248];
      88'b???????????????????????????????????????????????????????1????????????????????????????????:
        _14516_ = b[263:256];
      88'b??????????????????????????????????????????????????????1?????????????????????????????????:
        _14516_ = b[271:264];
      88'b?????????????????????????????????????????????????????1??????????????????????????????????:
        _14516_ = b[279:272];
      88'b????????????????????????????????????????????????????1???????????????????????????????????:
        _14516_ = b[287:280];
      88'b???????????????????????????????????????????????????1????????????????????????????????????:
        _14516_ = b[295:288];
      88'b??????????????????????????????????????????????????1?????????????????????????????????????:
        _14516_ = b[303:296];
      88'b?????????????????????????????????????????????????1??????????????????????????????????????:
        _14516_ = b[311:304];
      88'b????????????????????????????????????????????????1???????????????????????????????????????:
        _14516_ = b[319:312];
      88'b???????????????????????????????????????????????1????????????????????????????????????????:
        _14516_ = b[327:320];
      88'b??????????????????????????????????????????????1?????????????????????????????????????????:
        _14516_ = b[335:328];
      88'b?????????????????????????????????????????????1??????????????????????????????????????????:
        _14516_ = b[343:336];
      88'b????????????????????????????????????????????1???????????????????????????????????????????:
        _14516_ = b[351:344];
      88'b???????????????????????????????????????????1????????????????????????????????????????????:
        _14516_ = b[359:352];
      88'b??????????????????????????????????????????1?????????????????????????????????????????????:
        _14516_ = b[367:360];
      88'b?????????????????????????????????????????1??????????????????????????????????????????????:
        _14516_ = b[375:368];
      88'b????????????????????????????????????????1???????????????????????????????????????????????:
        _14516_ = b[383:376];
      88'b???????????????????????????????????????1????????????????????????????????????????????????:
        _14516_ = b[391:384];
      88'b??????????????????????????????????????1?????????????????????????????????????????????????:
        _14516_ = b[399:392];
      88'b?????????????????????????????????????1??????????????????????????????????????????????????:
        _14516_ = b[407:400];
      88'b????????????????????????????????????1???????????????????????????????????????????????????:
        _14516_ = b[415:408];
      88'b???????????????????????????????????1????????????????????????????????????????????????????:
        _14516_ = b[423:416];
      88'b??????????????????????????????????1?????????????????????????????????????????????????????:
        _14516_ = b[431:424];
      88'b?????????????????????????????????1??????????????????????????????????????????????????????:
        _14516_ = b[439:432];
      88'b????????????????????????????????1???????????????????????????????????????????????????????:
        _14516_ = b[447:440];
      88'b???????????????????????????????1????????????????????????????????????????????????????????:
        _14516_ = b[455:448];
      88'b??????????????????????????????1?????????????????????????????????????????????????????????:
        _14516_ = b[463:456];
      88'b?????????????????????????????1??????????????????????????????????????????????????????????:
        _14516_ = b[471:464];
      88'b????????????????????????????1???????????????????????????????????????????????????????????:
        _14516_ = b[479:472];
      88'b???????????????????????????1????????????????????????????????????????????????????????????:
        _14516_ = b[487:480];
      88'b??????????????????????????1?????????????????????????????????????????????????????????????:
        _14516_ = b[495:488];
      88'b?????????????????????????1??????????????????????????????????????????????????????????????:
        _14516_ = b[503:496];
      88'b????????????????????????1???????????????????????????????????????????????????????????????:
        _14516_ = b[511:504];
      88'b???????????????????????1????????????????????????????????????????????????????????????????:
        _14516_ = b[519:512];
      88'b??????????????????????1?????????????????????????????????????????????????????????????????:
        _14516_ = b[527:520];
      88'b?????????????????????1??????????????????????????????????????????????????????????????????:
        _14516_ = b[535:528];
      88'b????????????????????1???????????????????????????????????????????????????????????????????:
        _14516_ = b[543:536];
      88'b???????????????????1????????????????????????????????????????????????????????????????????:
        _14516_ = b[551:544];
      88'b??????????????????1?????????????????????????????????????????????????????????????????????:
        _14516_ = b[559:552];
      88'b?????????????????1??????????????????????????????????????????????????????????????????????:
        _14516_ = b[567:560];
      88'b????????????????1???????????????????????????????????????????????????????????????????????:
        _14516_ = b[575:568];
      88'b???????????????1????????????????????????????????????????????????????????????????????????:
        _14516_ = b[583:576];
      88'b??????????????1?????????????????????????????????????????????????????????????????????????:
        _14516_ = b[591:584];
      88'b?????????????1??????????????????????????????????????????????????????????????????????????:
        _14516_ = b[599:592];
      88'b????????????1???????????????????????????????????????????????????????????????????????????:
        _14516_ = b[607:600];
      88'b???????????1????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[615:608];
      88'b??????????1?????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[623:616];
      88'b?????????1??????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[631:624];
      88'b????????1???????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[639:632];
      88'b???????1????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[647:640];
      88'b??????1?????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[655:648];
      88'b?????1??????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[663:656];
      88'b????1???????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[671:664];
      88'b???1????????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[679:672];
      88'b??1?????????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[687:680];
      88'b?1??????????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[695:688];
      88'b1???????????????????????????????????????????????????????????????????????????????????????:
        _14516_ = b[703:696];
      default:
        _14516_ = a;
    endcase
  endfunction
  assign vec_data_087 = _14516_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688], data_d1[703:696] }, { _05173_, _05172_, _05171_, _05170_, _05169_, _05168_, _05167_, _05166_, _05165_, _05164_, _05163_, _05162_, _05161_, _05160_, _05159_, _05158_, _05157_, _05156_, _05155_, _05154_, _05153_, _05152_, _05151_, _05150_, _05149_, _05148_, _05147_, _05146_, _05145_, _05144_, _05143_, _05142_, _05141_, _05140_, _05139_, _05138_, _05137_, _05136_, _05135_, _05134_, _05133_, _05132_, _05131_, _05130_, _05129_, _05128_, _05127_, _05126_, _05125_, _05124_, _05123_, _05122_, _05121_, _05120_, _05119_, _05118_, _05117_, _05116_, _05115_, _05114_, _05113_, _05112_, _05111_, _05110_, _05109_, _05108_, _05107_, _05106_, _05105_, _05104_, _05103_, _05102_, _05101_, _05100_, _05099_, _05098_, _05097_, _05096_, _05095_, _05094_, _05093_, _05092_, _05091_, _05090_, _05089_, _05088_, _05087_, _05086_ });
  assign _05086_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1011000;
  assign _05087_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010111;
  assign _05088_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010110;
  assign _05089_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010101;
  assign _05090_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010100;
  assign _05091_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010011;
  assign _05092_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010010;
  assign _05093_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010001;
  assign _05094_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1010000;
  assign _05095_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001111;
  assign _05096_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001110;
  assign _05097_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001101;
  assign _05098_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001100;
  assign _05099_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001011;
  assign _05100_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001010;
  assign _05101_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001001;
  assign _05102_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1001000;
  assign _05103_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000111;
  assign _05104_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000110;
  assign _05105_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000101;
  assign _05106_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000100;
  assign _05107_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000011;
  assign _05108_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000010;
  assign _05109_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000001;
  assign _05110_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 7'b1000000;
  assign _05111_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111111;
  assign _05112_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111110;
  assign _05113_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111101;
  assign _05114_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111100;
  assign _05115_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111011;
  assign _05116_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111010;
  assign _05117_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111001;
  assign _05118_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b111000;
  assign _05119_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110111;
  assign _05120_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110110;
  assign _05121_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110101;
  assign _05122_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110100;
  assign _05123_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110011;
  assign _05124_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110010;
  assign _05125_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110001;
  assign _05126_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b110000;
  assign _05127_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101111;
  assign _05128_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101110;
  assign _05129_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101101;
  assign _05130_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101100;
  assign _05131_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101011;
  assign _05132_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101010;
  assign _05133_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101001;
  assign _05134_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b101000;
  assign _05135_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100111;
  assign _05136_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100110;
  assign _05137_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100101;
  assign _05138_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100100;
  assign _05139_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100011;
  assign _05140_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100010;
  assign _05141_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100001;
  assign _05142_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 6'b100000;
  assign _05143_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11111;
  assign _05144_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11110;
  assign _05145_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11101;
  assign _05146_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11100;
  assign _05147_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11011;
  assign _05148_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11010;
  assign _05149_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11001;
  assign _05150_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b11000;
  assign _05151_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10111;
  assign _05152_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10110;
  assign _05153_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10101;
  assign _05154_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10100;
  assign _05155_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10011;
  assign _05156_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10010;
  assign _05157_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10001;
  assign _05158_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 5'b10000;
  assign _05159_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1111;
  assign _05160_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1110;
  assign _05161_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1101;
  assign _05162_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1100;
  assign _05163_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1011;
  assign _05164_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1010;
  assign _05165_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1001;
  assign _05166_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 4'b1000;
  assign _05167_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 3'b111;
  assign _05168_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 3'b110;
  assign _05169_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 3'b101;
  assign _05170_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 3'b100;
  assign _05171_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 2'b11;
  assign _05172_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 2'b10;
  assign _05173_ = vec_sum_087_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8415" *) 1'b1;
  function [7:0] _14605_;
    input [7:0] a;
    input [695:0] b;
    input [86:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *)
    (* parallel_case *)
    casez (s)
      87'b??????????????????????????????????????????????????????????????????????????????????????1:
        _14605_ = b[7:0];
      87'b?????????????????????????????????????????????????????????????????????????????????????1?:
        _14605_ = b[15:8];
      87'b????????????????????????????????????????????????????????????????????????????????????1??:
        _14605_ = b[23:16];
      87'b???????????????????????????????????????????????????????????????????????????????????1???:
        _14605_ = b[31:24];
      87'b??????????????????????????????????????????????????????????????????????????????????1????:
        _14605_ = b[39:32];
      87'b?????????????????????????????????????????????????????????????????????????????????1?????:
        _14605_ = b[47:40];
      87'b????????????????????????????????????????????????????????????????????????????????1??????:
        _14605_ = b[55:48];
      87'b???????????????????????????????????????????????????????????????????????????????1???????:
        _14605_ = b[63:56];
      87'b??????????????????????????????????????????????????????????????????????????????1????????:
        _14605_ = b[71:64];
      87'b?????????????????????????????????????????????????????????????????????????????1?????????:
        _14605_ = b[79:72];
      87'b????????????????????????????????????????????????????????????????????????????1??????????:
        _14605_ = b[87:80];
      87'b???????????????????????????????????????????????????????????????????????????1???????????:
        _14605_ = b[95:88];
      87'b??????????????????????????????????????????????????????????????????????????1????????????:
        _14605_ = b[103:96];
      87'b?????????????????????????????????????????????????????????????????????????1?????????????:
        _14605_ = b[111:104];
      87'b????????????????????????????????????????????????????????????????????????1??????????????:
        _14605_ = b[119:112];
      87'b???????????????????????????????????????????????????????????????????????1???????????????:
        _14605_ = b[127:120];
      87'b??????????????????????????????????????????????????????????????????????1????????????????:
        _14605_ = b[135:128];
      87'b?????????????????????????????????????????????????????????????????????1?????????????????:
        _14605_ = b[143:136];
      87'b????????????????????????????????????????????????????????????????????1??????????????????:
        _14605_ = b[151:144];
      87'b???????????????????????????????????????????????????????????????????1???????????????????:
        _14605_ = b[159:152];
      87'b??????????????????????????????????????????????????????????????????1????????????????????:
        _14605_ = b[167:160];
      87'b?????????????????????????????????????????????????????????????????1?????????????????????:
        _14605_ = b[175:168];
      87'b????????????????????????????????????????????????????????????????1??????????????????????:
        _14605_ = b[183:176];
      87'b???????????????????????????????????????????????????????????????1???????????????????????:
        _14605_ = b[191:184];
      87'b??????????????????????????????????????????????????????????????1????????????????????????:
        _14605_ = b[199:192];
      87'b?????????????????????????????????????????????????????????????1?????????????????????????:
        _14605_ = b[207:200];
      87'b????????????????????????????????????????????????????????????1??????????????????????????:
        _14605_ = b[215:208];
      87'b???????????????????????????????????????????????????????????1???????????????????????????:
        _14605_ = b[223:216];
      87'b??????????????????????????????????????????????????????????1????????????????????????????:
        _14605_ = b[231:224];
      87'b?????????????????????????????????????????????????????????1?????????????????????????????:
        _14605_ = b[239:232];
      87'b????????????????????????????????????????????????????????1??????????????????????????????:
        _14605_ = b[247:240];
      87'b???????????????????????????????????????????????????????1???????????????????????????????:
        _14605_ = b[255:248];
      87'b??????????????????????????????????????????????????????1????????????????????????????????:
        _14605_ = b[263:256];
      87'b?????????????????????????????????????????????????????1?????????????????????????????????:
        _14605_ = b[271:264];
      87'b????????????????????????????????????????????????????1??????????????????????????????????:
        _14605_ = b[279:272];
      87'b???????????????????????????????????????????????????1???????????????????????????????????:
        _14605_ = b[287:280];
      87'b??????????????????????????????????????????????????1????????????????????????????????????:
        _14605_ = b[295:288];
      87'b?????????????????????????????????????????????????1?????????????????????????????????????:
        _14605_ = b[303:296];
      87'b????????????????????????????????????????????????1??????????????????????????????????????:
        _14605_ = b[311:304];
      87'b???????????????????????????????????????????????1???????????????????????????????????????:
        _14605_ = b[319:312];
      87'b??????????????????????????????????????????????1????????????????????????????????????????:
        _14605_ = b[327:320];
      87'b?????????????????????????????????????????????1?????????????????????????????????????????:
        _14605_ = b[335:328];
      87'b????????????????????????????????????????????1??????????????????????????????????????????:
        _14605_ = b[343:336];
      87'b???????????????????????????????????????????1???????????????????????????????????????????:
        _14605_ = b[351:344];
      87'b??????????????????????????????????????????1????????????????????????????????????????????:
        _14605_ = b[359:352];
      87'b?????????????????????????????????????????1?????????????????????????????????????????????:
        _14605_ = b[367:360];
      87'b????????????????????????????????????????1??????????????????????????????????????????????:
        _14605_ = b[375:368];
      87'b???????????????????????????????????????1???????????????????????????????????????????????:
        _14605_ = b[383:376];
      87'b??????????????????????????????????????1????????????????????????????????????????????????:
        _14605_ = b[391:384];
      87'b?????????????????????????????????????1?????????????????????????????????????????????????:
        _14605_ = b[399:392];
      87'b????????????????????????????????????1??????????????????????????????????????????????????:
        _14605_ = b[407:400];
      87'b???????????????????????????????????1???????????????????????????????????????????????????:
        _14605_ = b[415:408];
      87'b??????????????????????????????????1????????????????????????????????????????????????????:
        _14605_ = b[423:416];
      87'b?????????????????????????????????1?????????????????????????????????????????????????????:
        _14605_ = b[431:424];
      87'b????????????????????????????????1??????????????????????????????????????????????????????:
        _14605_ = b[439:432];
      87'b???????????????????????????????1???????????????????????????????????????????????????????:
        _14605_ = b[447:440];
      87'b??????????????????????????????1????????????????????????????????????????????????????????:
        _14605_ = b[455:448];
      87'b?????????????????????????????1?????????????????????????????????????????????????????????:
        _14605_ = b[463:456];
      87'b????????????????????????????1??????????????????????????????????????????????????????????:
        _14605_ = b[471:464];
      87'b???????????????????????????1???????????????????????????????????????????????????????????:
        _14605_ = b[479:472];
      87'b??????????????????????????1????????????????????????????????????????????????????????????:
        _14605_ = b[487:480];
      87'b?????????????????????????1?????????????????????????????????????????????????????????????:
        _14605_ = b[495:488];
      87'b????????????????????????1??????????????????????????????????????????????????????????????:
        _14605_ = b[503:496];
      87'b???????????????????????1???????????????????????????????????????????????????????????????:
        _14605_ = b[511:504];
      87'b??????????????????????1????????????????????????????????????????????????????????????????:
        _14605_ = b[519:512];
      87'b?????????????????????1?????????????????????????????????????????????????????????????????:
        _14605_ = b[527:520];
      87'b????????????????????1??????????????????????????????????????????????????????????????????:
        _14605_ = b[535:528];
      87'b???????????????????1???????????????????????????????????????????????????????????????????:
        _14605_ = b[543:536];
      87'b??????????????????1????????????????????????????????????????????????????????????????????:
        _14605_ = b[551:544];
      87'b?????????????????1?????????????????????????????????????????????????????????????????????:
        _14605_ = b[559:552];
      87'b????????????????1??????????????????????????????????????????????????????????????????????:
        _14605_ = b[567:560];
      87'b???????????????1???????????????????????????????????????????????????????????????????????:
        _14605_ = b[575:568];
      87'b??????????????1????????????????????????????????????????????????????????????????????????:
        _14605_ = b[583:576];
      87'b?????????????1?????????????????????????????????????????????????????????????????????????:
        _14605_ = b[591:584];
      87'b????????????1??????????????????????????????????????????????????????????????????????????:
        _14605_ = b[599:592];
      87'b???????????1???????????????????????????????????????????????????????????????????????????:
        _14605_ = b[607:600];
      87'b??????????1????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[615:608];
      87'b?????????1?????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[623:616];
      87'b????????1??????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[631:624];
      87'b???????1???????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[639:632];
      87'b??????1????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[647:640];
      87'b?????1?????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[655:648];
      87'b????1??????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[663:656];
      87'b???1???????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[671:664];
      87'b??1????????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[679:672];
      87'b?1?????????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[687:680];
      87'b1??????????????????????????????????????????????????????????????????????????????????????:
        _14605_ = b[695:688];
      default:
        _14605_ = a;
    endcase
  endfunction
  assign vec_data_086 = _14605_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680], data_d1[695:688] }, { _05260_, _05259_, _05258_, _05257_, _05256_, _05255_, _05254_, _05253_, _05252_, _05251_, _05250_, _05249_, _05248_, _05247_, _05246_, _05245_, _05244_, _05243_, _05242_, _05241_, _05240_, _05239_, _05238_, _05237_, _05236_, _05235_, _05234_, _05233_, _05232_, _05231_, _05230_, _05229_, _05228_, _05227_, _05226_, _05225_, _05224_, _05223_, _05222_, _05221_, _05220_, _05219_, _05218_, _05217_, _05216_, _05215_, _05214_, _05213_, _05212_, _05211_, _05210_, _05209_, _05208_, _05207_, _05206_, _05205_, _05204_, _05203_, _05202_, _05201_, _05200_, _05199_, _05198_, _05197_, _05196_, _05195_, _05194_, _05193_, _05192_, _05191_, _05190_, _05189_, _05188_, _05187_, _05186_, _05185_, _05184_, _05183_, _05182_, _05181_, _05180_, _05179_, _05178_, _05177_, _05176_, _05175_, _05174_ });
  assign _05174_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010111;
  assign _05175_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010110;
  assign _05176_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010101;
  assign _05177_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010100;
  assign _05178_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010011;
  assign _05179_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010010;
  assign _05180_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010001;
  assign _05181_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1010000;
  assign _05182_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001111;
  assign _05183_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001110;
  assign _05184_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001101;
  assign _05185_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001100;
  assign _05186_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001011;
  assign _05187_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001010;
  assign _05188_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001001;
  assign _05189_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1001000;
  assign _05190_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000111;
  assign _05191_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000110;
  assign _05192_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000101;
  assign _05193_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000100;
  assign _05194_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000011;
  assign _05195_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000010;
  assign _05196_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000001;
  assign _05197_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 7'b1000000;
  assign _05198_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111111;
  assign _05199_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111110;
  assign _05200_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111101;
  assign _05201_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111100;
  assign _05202_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111011;
  assign _05203_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111010;
  assign _05204_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111001;
  assign _05205_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b111000;
  assign _05206_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110111;
  assign _05207_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110110;
  assign _05208_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110101;
  assign _05209_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110100;
  assign _05210_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110011;
  assign _05211_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110010;
  assign _05212_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110001;
  assign _05213_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b110000;
  assign _05214_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101111;
  assign _05215_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101110;
  assign _05216_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101101;
  assign _05217_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101100;
  assign _05218_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101011;
  assign _05219_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101010;
  assign _05220_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101001;
  assign _05221_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b101000;
  assign _05222_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100111;
  assign _05223_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100110;
  assign _05224_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100101;
  assign _05225_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100100;
  assign _05226_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100011;
  assign _05227_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100010;
  assign _05228_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100001;
  assign _05229_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 6'b100000;
  assign _05230_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11111;
  assign _05231_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11110;
  assign _05232_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11101;
  assign _05233_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11100;
  assign _05234_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11011;
  assign _05235_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11010;
  assign _05236_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11001;
  assign _05237_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b11000;
  assign _05238_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10111;
  assign _05239_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10110;
  assign _05240_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10101;
  assign _05241_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10100;
  assign _05242_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10011;
  assign _05243_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10010;
  assign _05244_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10001;
  assign _05245_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 5'b10000;
  assign _05246_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1111;
  assign _05247_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1110;
  assign _05248_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1101;
  assign _05249_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1100;
  assign _05250_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1011;
  assign _05251_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1010;
  assign _05252_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1001;
  assign _05253_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 4'b1000;
  assign _05254_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 3'b111;
  assign _05255_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 3'b110;
  assign _05256_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 3'b101;
  assign _05257_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 3'b100;
  assign _05258_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 2'b11;
  assign _05259_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 2'b10;
  assign _05260_ = vec_sum_086_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8320" *) 1'b1;
  function [7:0] _14693_;
    input [7:0] a;
    input [687:0] b;
    input [85:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *)
    (* parallel_case *)
    casez (s)
      86'b?????????????????????????????????????????????????????????????????????????????????????1:
        _14693_ = b[7:0];
      86'b????????????????????????????????????????????????????????????????????????????????????1?:
        _14693_ = b[15:8];
      86'b???????????????????????????????????????????????????????????????????????????????????1??:
        _14693_ = b[23:16];
      86'b??????????????????????????????????????????????????????????????????????????????????1???:
        _14693_ = b[31:24];
      86'b?????????????????????????????????????????????????????????????????????????????????1????:
        _14693_ = b[39:32];
      86'b????????????????????????????????????????????????????????????????????????????????1?????:
        _14693_ = b[47:40];
      86'b???????????????????????????????????????????????????????????????????????????????1??????:
        _14693_ = b[55:48];
      86'b??????????????????????????????????????????????????????????????????????????????1???????:
        _14693_ = b[63:56];
      86'b?????????????????????????????????????????????????????????????????????????????1????????:
        _14693_ = b[71:64];
      86'b????????????????????????????????????????????????????????????????????????????1?????????:
        _14693_ = b[79:72];
      86'b???????????????????????????????????????????????????????????????????????????1??????????:
        _14693_ = b[87:80];
      86'b??????????????????????????????????????????????????????????????????????????1???????????:
        _14693_ = b[95:88];
      86'b?????????????????????????????????????????????????????????????????????????1????????????:
        _14693_ = b[103:96];
      86'b????????????????????????????????????????????????????????????????????????1?????????????:
        _14693_ = b[111:104];
      86'b???????????????????????????????????????????????????????????????????????1??????????????:
        _14693_ = b[119:112];
      86'b??????????????????????????????????????????????????????????????????????1???????????????:
        _14693_ = b[127:120];
      86'b?????????????????????????????????????????????????????????????????????1????????????????:
        _14693_ = b[135:128];
      86'b????????????????????????????????????????????????????????????????????1?????????????????:
        _14693_ = b[143:136];
      86'b???????????????????????????????????????????????????????????????????1??????????????????:
        _14693_ = b[151:144];
      86'b??????????????????????????????????????????????????????????????????1???????????????????:
        _14693_ = b[159:152];
      86'b?????????????????????????????????????????????????????????????????1????????????????????:
        _14693_ = b[167:160];
      86'b????????????????????????????????????????????????????????????????1?????????????????????:
        _14693_ = b[175:168];
      86'b???????????????????????????????????????????????????????????????1??????????????????????:
        _14693_ = b[183:176];
      86'b??????????????????????????????????????????????????????????????1???????????????????????:
        _14693_ = b[191:184];
      86'b?????????????????????????????????????????????????????????????1????????????????????????:
        _14693_ = b[199:192];
      86'b????????????????????????????????????????????????????????????1?????????????????????????:
        _14693_ = b[207:200];
      86'b???????????????????????????????????????????????????????????1??????????????????????????:
        _14693_ = b[215:208];
      86'b??????????????????????????????????????????????????????????1???????????????????????????:
        _14693_ = b[223:216];
      86'b?????????????????????????????????????????????????????????1????????????????????????????:
        _14693_ = b[231:224];
      86'b????????????????????????????????????????????????????????1?????????????????????????????:
        _14693_ = b[239:232];
      86'b???????????????????????????????????????????????????????1??????????????????????????????:
        _14693_ = b[247:240];
      86'b??????????????????????????????????????????????????????1???????????????????????????????:
        _14693_ = b[255:248];
      86'b?????????????????????????????????????????????????????1????????????????????????????????:
        _14693_ = b[263:256];
      86'b????????????????????????????????????????????????????1?????????????????????????????????:
        _14693_ = b[271:264];
      86'b???????????????????????????????????????????????????1??????????????????????????????????:
        _14693_ = b[279:272];
      86'b??????????????????????????????????????????????????1???????????????????????????????????:
        _14693_ = b[287:280];
      86'b?????????????????????????????????????????????????1????????????????????????????????????:
        _14693_ = b[295:288];
      86'b????????????????????????????????????????????????1?????????????????????????????????????:
        _14693_ = b[303:296];
      86'b???????????????????????????????????????????????1??????????????????????????????????????:
        _14693_ = b[311:304];
      86'b??????????????????????????????????????????????1???????????????????????????????????????:
        _14693_ = b[319:312];
      86'b?????????????????????????????????????????????1????????????????????????????????????????:
        _14693_ = b[327:320];
      86'b????????????????????????????????????????????1?????????????????????????????????????????:
        _14693_ = b[335:328];
      86'b???????????????????????????????????????????1??????????????????????????????????????????:
        _14693_ = b[343:336];
      86'b??????????????????????????????????????????1???????????????????????????????????????????:
        _14693_ = b[351:344];
      86'b?????????????????????????????????????????1????????????????????????????????????????????:
        _14693_ = b[359:352];
      86'b????????????????????????????????????????1?????????????????????????????????????????????:
        _14693_ = b[367:360];
      86'b???????????????????????????????????????1??????????????????????????????????????????????:
        _14693_ = b[375:368];
      86'b??????????????????????????????????????1???????????????????????????????????????????????:
        _14693_ = b[383:376];
      86'b?????????????????????????????????????1????????????????????????????????????????????????:
        _14693_ = b[391:384];
      86'b????????????????????????????????????1?????????????????????????????????????????????????:
        _14693_ = b[399:392];
      86'b???????????????????????????????????1??????????????????????????????????????????????????:
        _14693_ = b[407:400];
      86'b??????????????????????????????????1???????????????????????????????????????????????????:
        _14693_ = b[415:408];
      86'b?????????????????????????????????1????????????????????????????????????????????????????:
        _14693_ = b[423:416];
      86'b????????????????????????????????1?????????????????????????????????????????????????????:
        _14693_ = b[431:424];
      86'b???????????????????????????????1??????????????????????????????????????????????????????:
        _14693_ = b[439:432];
      86'b??????????????????????????????1???????????????????????????????????????????????????????:
        _14693_ = b[447:440];
      86'b?????????????????????????????1????????????????????????????????????????????????????????:
        _14693_ = b[455:448];
      86'b????????????????????????????1?????????????????????????????????????????????????????????:
        _14693_ = b[463:456];
      86'b???????????????????????????1??????????????????????????????????????????????????????????:
        _14693_ = b[471:464];
      86'b??????????????????????????1???????????????????????????????????????????????????????????:
        _14693_ = b[479:472];
      86'b?????????????????????????1????????????????????????????????????????????????????????????:
        _14693_ = b[487:480];
      86'b????????????????????????1?????????????????????????????????????????????????????????????:
        _14693_ = b[495:488];
      86'b???????????????????????1??????????????????????????????????????????????????????????????:
        _14693_ = b[503:496];
      86'b??????????????????????1???????????????????????????????????????????????????????????????:
        _14693_ = b[511:504];
      86'b?????????????????????1????????????????????????????????????????????????????????????????:
        _14693_ = b[519:512];
      86'b????????????????????1?????????????????????????????????????????????????????????????????:
        _14693_ = b[527:520];
      86'b???????????????????1??????????????????????????????????????????????????????????????????:
        _14693_ = b[535:528];
      86'b??????????????????1???????????????????????????????????????????????????????????????????:
        _14693_ = b[543:536];
      86'b?????????????????1????????????????????????????????????????????????????????????????????:
        _14693_ = b[551:544];
      86'b????????????????1?????????????????????????????????????????????????????????????????????:
        _14693_ = b[559:552];
      86'b???????????????1??????????????????????????????????????????????????????????????????????:
        _14693_ = b[567:560];
      86'b??????????????1???????????????????????????????????????????????????????????????????????:
        _14693_ = b[575:568];
      86'b?????????????1????????????????????????????????????????????????????????????????????????:
        _14693_ = b[583:576];
      86'b????????????1?????????????????????????????????????????????????????????????????????????:
        _14693_ = b[591:584];
      86'b???????????1??????????????????????????????????????????????????????????????????????????:
        _14693_ = b[599:592];
      86'b??????????1???????????????????????????????????????????????????????????????????????????:
        _14693_ = b[607:600];
      86'b?????????1????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[615:608];
      86'b????????1?????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[623:616];
      86'b???????1??????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[631:624];
      86'b??????1???????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[639:632];
      86'b?????1????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[647:640];
      86'b????1?????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[655:648];
      86'b???1??????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[663:656];
      86'b??1???????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[671:664];
      86'b?1????????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[679:672];
      86'b1?????????????????????????????????????????????????????????????????????????????????????:
        _14693_ = b[687:680];
      default:
        _14693_ = a;
    endcase
  endfunction
  assign vec_data_085 = _14693_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672], data_d1[687:680] }, { _05346_, _05345_, _05344_, _05343_, _05342_, _05341_, _05340_, _05339_, _05338_, _05337_, _05336_, _05335_, _05334_, _05333_, _05332_, _05331_, _05330_, _05329_, _05328_, _05327_, _05326_, _05325_, _05324_, _05323_, _05322_, _05321_, _05320_, _05319_, _05318_, _05317_, _05316_, _05315_, _05314_, _05313_, _05312_, _05311_, _05310_, _05309_, _05308_, _05307_, _05306_, _05305_, _05304_, _05303_, _05302_, _05301_, _05300_, _05299_, _05298_, _05297_, _05296_, _05295_, _05294_, _05293_, _05292_, _05291_, _05290_, _05289_, _05288_, _05287_, _05286_, _05285_, _05284_, _05283_, _05282_, _05281_, _05280_, _05279_, _05278_, _05277_, _05276_, _05275_, _05274_, _05273_, _05272_, _05271_, _05270_, _05269_, _05268_, _05267_, _05266_, _05265_, _05264_, _05263_, _05262_, _05261_ });
  assign _05261_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010110;
  assign _05262_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010101;
  assign _05263_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010100;
  assign _05264_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010011;
  assign _05265_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010010;
  assign _05266_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010001;
  assign _05267_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1010000;
  assign _05268_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001111;
  assign _05269_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001110;
  assign _05270_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001101;
  assign _05271_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001100;
  assign _05272_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001011;
  assign _05273_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001010;
  assign _05274_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001001;
  assign _05275_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1001000;
  assign _05276_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000111;
  assign _05277_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000110;
  assign _05278_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000101;
  assign _05279_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000100;
  assign _05280_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000011;
  assign _05281_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000010;
  assign _05282_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000001;
  assign _05283_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 7'b1000000;
  assign _05284_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111111;
  assign _05285_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111110;
  assign _05286_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111101;
  assign _05287_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111100;
  assign _05288_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111011;
  assign _05289_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111010;
  assign _05290_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111001;
  assign _05291_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b111000;
  assign _05292_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110111;
  assign _05293_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110110;
  assign _05294_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110101;
  assign _05295_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110100;
  assign _05296_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110011;
  assign _05297_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110010;
  assign _05298_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110001;
  assign _05299_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b110000;
  assign _05300_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101111;
  assign _05301_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101110;
  assign _05302_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101101;
  assign _05303_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101100;
  assign _05304_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101011;
  assign _05305_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101010;
  assign _05306_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101001;
  assign _05307_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b101000;
  assign _05308_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100111;
  assign _05309_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100110;
  assign _05310_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100101;
  assign _05311_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100100;
  assign _05312_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100011;
  assign _05313_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100010;
  assign _05314_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100001;
  assign _05315_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 6'b100000;
  assign _05316_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11111;
  assign _05317_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11110;
  assign _05318_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11101;
  assign _05319_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11100;
  assign _05320_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11011;
  assign _05321_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11010;
  assign _05322_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11001;
  assign _05323_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b11000;
  assign _05324_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10111;
  assign _05325_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10110;
  assign _05326_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10101;
  assign _05327_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10100;
  assign _05328_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10011;
  assign _05329_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10010;
  assign _05330_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10001;
  assign _05331_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 5'b10000;
  assign _05332_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1111;
  assign _05333_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1110;
  assign _05334_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1101;
  assign _05335_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1100;
  assign _05336_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1011;
  assign _05337_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1010;
  assign _05338_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1001;
  assign _05339_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 4'b1000;
  assign _05340_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8233|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 3'b111;
  assign _05341_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 3'b110;
  assign _05342_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 3'b101;
  assign _05343_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 3'b100;
  assign _05344_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 2'b11;
  assign _05345_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 2'b10;
  assign _05346_ = vec_sum_085_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8226" *) 1'b1;
  function [7:0] _14780_;
    input [7:0] a;
    input [679:0] b;
    input [84:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *)
    (* parallel_case *)
    casez (s)
      85'b????????????????????????????????????????????????????????????????????????????????????1:
        _14780_ = b[7:0];
      85'b???????????????????????????????????????????????????????????????????????????????????1?:
        _14780_ = b[15:8];
      85'b??????????????????????????????????????????????????????????????????????????????????1??:
        _14780_ = b[23:16];
      85'b?????????????????????????????????????????????????????????????????????????????????1???:
        _14780_ = b[31:24];
      85'b????????????????????????????????????????????????????????????????????????????????1????:
        _14780_ = b[39:32];
      85'b???????????????????????????????????????????????????????????????????????????????1?????:
        _14780_ = b[47:40];
      85'b??????????????????????????????????????????????????????????????????????????????1??????:
        _14780_ = b[55:48];
      85'b?????????????????????????????????????????????????????????????????????????????1???????:
        _14780_ = b[63:56];
      85'b????????????????????????????????????????????????????????????????????????????1????????:
        _14780_ = b[71:64];
      85'b???????????????????????????????????????????????????????????????????????????1?????????:
        _14780_ = b[79:72];
      85'b??????????????????????????????????????????????????????????????????????????1??????????:
        _14780_ = b[87:80];
      85'b?????????????????????????????????????????????????????????????????????????1???????????:
        _14780_ = b[95:88];
      85'b????????????????????????????????????????????????????????????????????????1????????????:
        _14780_ = b[103:96];
      85'b???????????????????????????????????????????????????????????????????????1?????????????:
        _14780_ = b[111:104];
      85'b??????????????????????????????????????????????????????????????????????1??????????????:
        _14780_ = b[119:112];
      85'b?????????????????????????????????????????????????????????????????????1???????????????:
        _14780_ = b[127:120];
      85'b????????????????????????????????????????????????????????????????????1????????????????:
        _14780_ = b[135:128];
      85'b???????????????????????????????????????????????????????????????????1?????????????????:
        _14780_ = b[143:136];
      85'b??????????????????????????????????????????????????????????????????1??????????????????:
        _14780_ = b[151:144];
      85'b?????????????????????????????????????????????????????????????????1???????????????????:
        _14780_ = b[159:152];
      85'b????????????????????????????????????????????????????????????????1????????????????????:
        _14780_ = b[167:160];
      85'b???????????????????????????????????????????????????????????????1?????????????????????:
        _14780_ = b[175:168];
      85'b??????????????????????????????????????????????????????????????1??????????????????????:
        _14780_ = b[183:176];
      85'b?????????????????????????????????????????????????????????????1???????????????????????:
        _14780_ = b[191:184];
      85'b????????????????????????????????????????????????????????????1????????????????????????:
        _14780_ = b[199:192];
      85'b???????????????????????????????????????????????????????????1?????????????????????????:
        _14780_ = b[207:200];
      85'b??????????????????????????????????????????????????????????1??????????????????????????:
        _14780_ = b[215:208];
      85'b?????????????????????????????????????????????????????????1???????????????????????????:
        _14780_ = b[223:216];
      85'b????????????????????????????????????????????????????????1????????????????????????????:
        _14780_ = b[231:224];
      85'b???????????????????????????????????????????????????????1?????????????????????????????:
        _14780_ = b[239:232];
      85'b??????????????????????????????????????????????????????1??????????????????????????????:
        _14780_ = b[247:240];
      85'b?????????????????????????????????????????????????????1???????????????????????????????:
        _14780_ = b[255:248];
      85'b????????????????????????????????????????????????????1????????????????????????????????:
        _14780_ = b[263:256];
      85'b???????????????????????????????????????????????????1?????????????????????????????????:
        _14780_ = b[271:264];
      85'b??????????????????????????????????????????????????1??????????????????????????????????:
        _14780_ = b[279:272];
      85'b?????????????????????????????????????????????????1???????????????????????????????????:
        _14780_ = b[287:280];
      85'b????????????????????????????????????????????????1????????????????????????????????????:
        _14780_ = b[295:288];
      85'b???????????????????????????????????????????????1?????????????????????????????????????:
        _14780_ = b[303:296];
      85'b??????????????????????????????????????????????1??????????????????????????????????????:
        _14780_ = b[311:304];
      85'b?????????????????????????????????????????????1???????????????????????????????????????:
        _14780_ = b[319:312];
      85'b????????????????????????????????????????????1????????????????????????????????????????:
        _14780_ = b[327:320];
      85'b???????????????????????????????????????????1?????????????????????????????????????????:
        _14780_ = b[335:328];
      85'b??????????????????????????????????????????1??????????????????????????????????????????:
        _14780_ = b[343:336];
      85'b?????????????????????????????????????????1???????????????????????????????????????????:
        _14780_ = b[351:344];
      85'b????????????????????????????????????????1????????????????????????????????????????????:
        _14780_ = b[359:352];
      85'b???????????????????????????????????????1?????????????????????????????????????????????:
        _14780_ = b[367:360];
      85'b??????????????????????????????????????1??????????????????????????????????????????????:
        _14780_ = b[375:368];
      85'b?????????????????????????????????????1???????????????????????????????????????????????:
        _14780_ = b[383:376];
      85'b????????????????????????????????????1????????????????????????????????????????????????:
        _14780_ = b[391:384];
      85'b???????????????????????????????????1?????????????????????????????????????????????????:
        _14780_ = b[399:392];
      85'b??????????????????????????????????1??????????????????????????????????????????????????:
        _14780_ = b[407:400];
      85'b?????????????????????????????????1???????????????????????????????????????????????????:
        _14780_ = b[415:408];
      85'b????????????????????????????????1????????????????????????????????????????????????????:
        _14780_ = b[423:416];
      85'b???????????????????????????????1?????????????????????????????????????????????????????:
        _14780_ = b[431:424];
      85'b??????????????????????????????1??????????????????????????????????????????????????????:
        _14780_ = b[439:432];
      85'b?????????????????????????????1???????????????????????????????????????????????????????:
        _14780_ = b[447:440];
      85'b????????????????????????????1????????????????????????????????????????????????????????:
        _14780_ = b[455:448];
      85'b???????????????????????????1?????????????????????????????????????????????????????????:
        _14780_ = b[463:456];
      85'b??????????????????????????1??????????????????????????????????????????????????????????:
        _14780_ = b[471:464];
      85'b?????????????????????????1???????????????????????????????????????????????????????????:
        _14780_ = b[479:472];
      85'b????????????????????????1????????????????????????????????????????????????????????????:
        _14780_ = b[487:480];
      85'b???????????????????????1?????????????????????????????????????????????????????????????:
        _14780_ = b[495:488];
      85'b??????????????????????1??????????????????????????????????????????????????????????????:
        _14780_ = b[503:496];
      85'b?????????????????????1???????????????????????????????????????????????????????????????:
        _14780_ = b[511:504];
      85'b????????????????????1????????????????????????????????????????????????????????????????:
        _14780_ = b[519:512];
      85'b???????????????????1?????????????????????????????????????????????????????????????????:
        _14780_ = b[527:520];
      85'b??????????????????1??????????????????????????????????????????????????????????????????:
        _14780_ = b[535:528];
      85'b?????????????????1???????????????????????????????????????????????????????????????????:
        _14780_ = b[543:536];
      85'b????????????????1????????????????????????????????????????????????????????????????????:
        _14780_ = b[551:544];
      85'b???????????????1?????????????????????????????????????????????????????????????????????:
        _14780_ = b[559:552];
      85'b??????????????1??????????????????????????????????????????????????????????????????????:
        _14780_ = b[567:560];
      85'b?????????????1???????????????????????????????????????????????????????????????????????:
        _14780_ = b[575:568];
      85'b????????????1????????????????????????????????????????????????????????????????????????:
        _14780_ = b[583:576];
      85'b???????????1?????????????????????????????????????????????????????????????????????????:
        _14780_ = b[591:584];
      85'b??????????1??????????????????????????????????????????????????????????????????????????:
        _14780_ = b[599:592];
      85'b?????????1???????????????????????????????????????????????????????????????????????????:
        _14780_ = b[607:600];
      85'b????????1????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[615:608];
      85'b???????1?????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[623:616];
      85'b??????1??????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[631:624];
      85'b?????1???????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[639:632];
      85'b????1????????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[647:640];
      85'b???1?????????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[655:648];
      85'b??1??????????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[663:656];
      85'b?1???????????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[671:664];
      85'b1????????????????????????????????????????????????????????????????????????????????????:
        _14780_ = b[679:672];
      default:
        _14780_ = a;
    endcase
  endfunction
  assign vec_data_084 = _14780_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664], data_d1[679:672] }, { _05431_, _05430_, _05429_, _05428_, _05427_, _05426_, _05425_, _05424_, _05423_, _05422_, _05421_, _05420_, _05419_, _05418_, _05417_, _05416_, _05415_, _05414_, _05413_, _05412_, _05411_, _05410_, _05409_, _05408_, _05407_, _05406_, _05405_, _05404_, _05403_, _05402_, _05401_, _05400_, _05399_, _05398_, _05397_, _05396_, _05395_, _05394_, _05393_, _05392_, _05391_, _05390_, _05389_, _05388_, _05387_, _05386_, _05385_, _05384_, _05383_, _05382_, _05381_, _05380_, _05379_, _05378_, _05377_, _05376_, _05375_, _05374_, _05373_, _05372_, _05371_, _05370_, _05369_, _05368_, _05367_, _05366_, _05365_, _05364_, _05363_, _05362_, _05361_, _05360_, _05359_, _05358_, _05357_, _05356_, _05355_, _05354_, _05353_, _05352_, _05351_, _05350_, _05349_, _05348_, _05347_ });
  assign _05347_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010101;
  assign _05348_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010100;
  assign _05349_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010011;
  assign _05350_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010010;
  assign _05351_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010001;
  assign _05352_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1010000;
  assign _05353_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001111;
  assign _05354_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001110;
  assign _05355_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001101;
  assign _05356_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001100;
  assign _05357_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001011;
  assign _05358_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001010;
  assign _05359_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001001;
  assign _05360_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1001000;
  assign _05361_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000111;
  assign _05362_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000110;
  assign _05363_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000101;
  assign _05364_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000100;
  assign _05365_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000011;
  assign _05366_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000010;
  assign _05367_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000001;
  assign _05368_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 7'b1000000;
  assign _05369_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111111;
  assign _05370_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111110;
  assign _05371_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111101;
  assign _05372_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111100;
  assign _05373_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111011;
  assign _05374_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111010;
  assign _05375_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111001;
  assign _05376_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b111000;
  assign _05377_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110111;
  assign _05378_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110110;
  assign _05379_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110101;
  assign _05380_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110100;
  assign _05381_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110011;
  assign _05382_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110010;
  assign _05383_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110001;
  assign _05384_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b110000;
  assign _05385_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101111;
  assign _05386_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101110;
  assign _05387_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101101;
  assign _05388_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101100;
  assign _05389_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8176|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101011;
  assign _05390_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101010;
  assign _05391_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101001;
  assign _05392_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b101000;
  assign _05393_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100111;
  assign _05394_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100110;
  assign _05395_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100101;
  assign _05396_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100100;
  assign _05397_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100011;
  assign _05398_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100010;
  assign _05399_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100001;
  assign _05400_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 6'b100000;
  assign _05401_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11111;
  assign _05402_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11110;
  assign _05403_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11101;
  assign _05404_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11100;
  assign _05405_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11011;
  assign _05406_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11010;
  assign _05407_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11001;
  assign _05408_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b11000;
  assign _05409_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10111;
  assign _05410_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10110;
  assign _05411_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10101;
  assign _05412_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10100;
  assign _05413_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10011;
  assign _05414_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10010;
  assign _05415_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10001;
  assign _05416_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 5'b10000;
  assign _05417_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1111;
  assign _05418_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1110;
  assign _05419_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1101;
  assign _05420_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1100;
  assign _05421_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1011;
  assign _05422_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1010;
  assign _05423_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1001;
  assign _05424_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 4'b1000;
  assign _05425_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 3'b111;
  assign _05426_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 3'b110;
  assign _05427_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 3'b101;
  assign _05428_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 3'b100;
  assign _05429_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 2'b11;
  assign _05430_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 2'b10;
  assign _05431_ = vec_sum_084_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8133" *) 1'b1;
  function [7:0] _14866_;
    input [7:0] a;
    input [671:0] b;
    input [83:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *)
    (* parallel_case *)
    casez (s)
      84'b???????????????????????????????????????????????????????????????????????????????????1:
        _14866_ = b[7:0];
      84'b??????????????????????????????????????????????????????????????????????????????????1?:
        _14866_ = b[15:8];
      84'b?????????????????????????????????????????????????????????????????????????????????1??:
        _14866_ = b[23:16];
      84'b????????????????????????????????????????????????????????????????????????????????1???:
        _14866_ = b[31:24];
      84'b???????????????????????????????????????????????????????????????????????????????1????:
        _14866_ = b[39:32];
      84'b??????????????????????????????????????????????????????????????????????????????1?????:
        _14866_ = b[47:40];
      84'b?????????????????????????????????????????????????????????????????????????????1??????:
        _14866_ = b[55:48];
      84'b????????????????????????????????????????????????????????????????????????????1???????:
        _14866_ = b[63:56];
      84'b???????????????????????????????????????????????????????????????????????????1????????:
        _14866_ = b[71:64];
      84'b??????????????????????????????????????????????????????????????????????????1?????????:
        _14866_ = b[79:72];
      84'b?????????????????????????????????????????????????????????????????????????1??????????:
        _14866_ = b[87:80];
      84'b????????????????????????????????????????????????????????????????????????1???????????:
        _14866_ = b[95:88];
      84'b???????????????????????????????????????????????????????????????????????1????????????:
        _14866_ = b[103:96];
      84'b??????????????????????????????????????????????????????????????????????1?????????????:
        _14866_ = b[111:104];
      84'b?????????????????????????????????????????????????????????????????????1??????????????:
        _14866_ = b[119:112];
      84'b????????????????????????????????????????????????????????????????????1???????????????:
        _14866_ = b[127:120];
      84'b???????????????????????????????????????????????????????????????????1????????????????:
        _14866_ = b[135:128];
      84'b??????????????????????????????????????????????????????????????????1?????????????????:
        _14866_ = b[143:136];
      84'b?????????????????????????????????????????????????????????????????1??????????????????:
        _14866_ = b[151:144];
      84'b????????????????????????????????????????????????????????????????1???????????????????:
        _14866_ = b[159:152];
      84'b???????????????????????????????????????????????????????????????1????????????????????:
        _14866_ = b[167:160];
      84'b??????????????????????????????????????????????????????????????1?????????????????????:
        _14866_ = b[175:168];
      84'b?????????????????????????????????????????????????????????????1??????????????????????:
        _14866_ = b[183:176];
      84'b????????????????????????????????????????????????????????????1???????????????????????:
        _14866_ = b[191:184];
      84'b???????????????????????????????????????????????????????????1????????????????????????:
        _14866_ = b[199:192];
      84'b??????????????????????????????????????????????????????????1?????????????????????????:
        _14866_ = b[207:200];
      84'b?????????????????????????????????????????????????????????1??????????????????????????:
        _14866_ = b[215:208];
      84'b????????????????????????????????????????????????????????1???????????????????????????:
        _14866_ = b[223:216];
      84'b???????????????????????????????????????????????????????1????????????????????????????:
        _14866_ = b[231:224];
      84'b??????????????????????????????????????????????????????1?????????????????????????????:
        _14866_ = b[239:232];
      84'b?????????????????????????????????????????????????????1??????????????????????????????:
        _14866_ = b[247:240];
      84'b????????????????????????????????????????????????????1???????????????????????????????:
        _14866_ = b[255:248];
      84'b???????????????????????????????????????????????????1????????????????????????????????:
        _14866_ = b[263:256];
      84'b??????????????????????????????????????????????????1?????????????????????????????????:
        _14866_ = b[271:264];
      84'b?????????????????????????????????????????????????1??????????????????????????????????:
        _14866_ = b[279:272];
      84'b????????????????????????????????????????????????1???????????????????????????????????:
        _14866_ = b[287:280];
      84'b???????????????????????????????????????????????1????????????????????????????????????:
        _14866_ = b[295:288];
      84'b??????????????????????????????????????????????1?????????????????????????????????????:
        _14866_ = b[303:296];
      84'b?????????????????????????????????????????????1??????????????????????????????????????:
        _14866_ = b[311:304];
      84'b????????????????????????????????????????????1???????????????????????????????????????:
        _14866_ = b[319:312];
      84'b???????????????????????????????????????????1????????????????????????????????????????:
        _14866_ = b[327:320];
      84'b??????????????????????????????????????????1?????????????????????????????????????????:
        _14866_ = b[335:328];
      84'b?????????????????????????????????????????1??????????????????????????????????????????:
        _14866_ = b[343:336];
      84'b????????????????????????????????????????1???????????????????????????????????????????:
        _14866_ = b[351:344];
      84'b???????????????????????????????????????1????????????????????????????????????????????:
        _14866_ = b[359:352];
      84'b??????????????????????????????????????1?????????????????????????????????????????????:
        _14866_ = b[367:360];
      84'b?????????????????????????????????????1??????????????????????????????????????????????:
        _14866_ = b[375:368];
      84'b????????????????????????????????????1???????????????????????????????????????????????:
        _14866_ = b[383:376];
      84'b???????????????????????????????????1????????????????????????????????????????????????:
        _14866_ = b[391:384];
      84'b??????????????????????????????????1?????????????????????????????????????????????????:
        _14866_ = b[399:392];
      84'b?????????????????????????????????1??????????????????????????????????????????????????:
        _14866_ = b[407:400];
      84'b????????????????????????????????1???????????????????????????????????????????????????:
        _14866_ = b[415:408];
      84'b???????????????????????????????1????????????????????????????????????????????????????:
        _14866_ = b[423:416];
      84'b??????????????????????????????1?????????????????????????????????????????????????????:
        _14866_ = b[431:424];
      84'b?????????????????????????????1??????????????????????????????????????????????????????:
        _14866_ = b[439:432];
      84'b????????????????????????????1???????????????????????????????????????????????????????:
        _14866_ = b[447:440];
      84'b???????????????????????????1????????????????????????????????????????????????????????:
        _14866_ = b[455:448];
      84'b??????????????????????????1?????????????????????????????????????????????????????????:
        _14866_ = b[463:456];
      84'b?????????????????????????1??????????????????????????????????????????????????????????:
        _14866_ = b[471:464];
      84'b????????????????????????1???????????????????????????????????????????????????????????:
        _14866_ = b[479:472];
      84'b???????????????????????1????????????????????????????????????????????????????????????:
        _14866_ = b[487:480];
      84'b??????????????????????1?????????????????????????????????????????????????????????????:
        _14866_ = b[495:488];
      84'b?????????????????????1??????????????????????????????????????????????????????????????:
        _14866_ = b[503:496];
      84'b????????????????????1???????????????????????????????????????????????????????????????:
        _14866_ = b[511:504];
      84'b???????????????????1????????????????????????????????????????????????????????????????:
        _14866_ = b[519:512];
      84'b??????????????????1?????????????????????????????????????????????????????????????????:
        _14866_ = b[527:520];
      84'b?????????????????1??????????????????????????????????????????????????????????????????:
        _14866_ = b[535:528];
      84'b????????????????1???????????????????????????????????????????????????????????????????:
        _14866_ = b[543:536];
      84'b???????????????1????????????????????????????????????????????????????????????????????:
        _14866_ = b[551:544];
      84'b??????????????1?????????????????????????????????????????????????????????????????????:
        _14866_ = b[559:552];
      84'b?????????????1??????????????????????????????????????????????????????????????????????:
        _14866_ = b[567:560];
      84'b????????????1???????????????????????????????????????????????????????????????????????:
        _14866_ = b[575:568];
      84'b???????????1????????????????????????????????????????????????????????????????????????:
        _14866_ = b[583:576];
      84'b??????????1?????????????????????????????????????????????????????????????????????????:
        _14866_ = b[591:584];
      84'b?????????1??????????????????????????????????????????????????????????????????????????:
        _14866_ = b[599:592];
      84'b????????1???????????????????????????????????????????????????????????????????????????:
        _14866_ = b[607:600];
      84'b???????1????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[615:608];
      84'b??????1?????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[623:616];
      84'b?????1??????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[631:624];
      84'b????1???????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[639:632];
      84'b???1????????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[647:640];
      84'b??1?????????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[655:648];
      84'b?1??????????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[663:656];
      84'b1???????????????????????????????????????????????????????????????????????????????????:
        _14866_ = b[671:664];
      default:
        _14866_ = a;
    endcase
  endfunction
  assign vec_data_083 = _14866_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656], data_d1[671:664] }, { _05515_, _05514_, _05513_, _05512_, _05511_, _05510_, _05509_, _05508_, _05507_, _05506_, _05505_, _05504_, _05503_, _05502_, _05501_, _05500_, _05499_, _05498_, _05497_, _05496_, _05495_, _05494_, _05493_, _05492_, _05491_, _05490_, _05489_, _05488_, _05487_, _05486_, _05485_, _05484_, _05483_, _05482_, _05481_, _05480_, _05479_, _05478_, _05477_, _05476_, _05475_, _05474_, _05473_, _05472_, _05471_, _05470_, _05469_, _05468_, _05467_, _05466_, _05465_, _05464_, _05463_, _05462_, _05461_, _05460_, _05459_, _05458_, _05457_, _05456_, _05455_, _05454_, _05453_, _05452_, _05451_, _05450_, _05449_, _05448_, _05447_, _05446_, _05445_, _05444_, _05443_, _05442_, _05441_, _05440_, _05439_, _05438_, _05437_, _05436_, _05435_, _05434_, _05433_, _05432_ });
  assign _05432_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1010100;
  assign _05433_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1010011;
  assign _05434_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1010010;
  assign _05435_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1010001;
  assign _05436_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1010000;
  assign _05437_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001111;
  assign _05438_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001110;
  assign _05439_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001101;
  assign _05440_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001100;
  assign _05441_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001011;
  assign _05442_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001010;
  assign _05443_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001001;
  assign _05444_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1001000;
  assign _05445_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000111;
  assign _05446_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000110;
  assign _05447_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000101;
  assign _05448_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000100;
  assign _05449_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000011;
  assign _05450_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000010;
  assign _05451_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000001;
  assign _05452_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 7'b1000000;
  assign _05453_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111111;
  assign _05454_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111110;
  assign _05455_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111101;
  assign _05456_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111100;
  assign _05457_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111011;
  assign _05458_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111010;
  assign _05459_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111001;
  assign _05460_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b111000;
  assign _05461_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110111;
  assign _05462_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110110;
  assign _05463_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110101;
  assign _05464_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110100;
  assign _05465_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110011;
  assign _05466_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110010;
  assign _05467_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110001;
  assign _05468_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b110000;
  assign _05469_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101111;
  assign _05470_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101110;
  assign _05471_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101101;
  assign _05472_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101100;
  assign _05473_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101011;
  assign _05474_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101010;
  assign _05475_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101001;
  assign _05476_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b101000;
  assign _05477_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100111;
  assign _05478_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100110;
  assign _05479_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100101;
  assign _05480_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100100;
  assign _05481_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100011;
  assign _05482_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100010;
  assign _05483_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100001;
  assign _05484_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 6'b100000;
  assign _05485_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11111;
  assign _05486_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11110;
  assign _05487_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11101;
  assign _05488_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11100;
  assign _05489_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11011;
  assign _05490_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11010;
  assign _05491_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11001;
  assign _05492_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b11000;
  assign _05493_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10111;
  assign _05494_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10110;
  assign _05495_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10101;
  assign _05496_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10100;
  assign _05497_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10011;
  assign _05498_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10010;
  assign _05499_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10001;
  assign _05500_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 5'b10000;
  assign _05501_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1111;
  assign _05502_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1110;
  assign _05503_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1101;
  assign _05504_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1100;
  assign _05505_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1011;
  assign _05506_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1010;
  assign _05507_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1001;
  assign _05508_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 4'b1000;
  assign _05509_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 3'b111;
  assign _05510_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 3'b110;
  assign _05511_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 3'b101;
  assign _05512_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 3'b100;
  assign _05513_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 2'b11;
  assign _05514_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 2'b10;
  assign _05515_ = vec_sum_083_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8041" *) 1'b1;
  function [7:0] _14951_;
    input [7:0] a;
    input [663:0] b;
    input [82:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *)
    (* parallel_case *)
    casez (s)
      83'b??????????????????????????????????????????????????????????????????????????????????1:
        _14951_ = b[7:0];
      83'b?????????????????????????????????????????????????????????????????????????????????1?:
        _14951_ = b[15:8];
      83'b????????????????????????????????????????????????????????????????????????????????1??:
        _14951_ = b[23:16];
      83'b???????????????????????????????????????????????????????????????????????????????1???:
        _14951_ = b[31:24];
      83'b??????????????????????????????????????????????????????????????????????????????1????:
        _14951_ = b[39:32];
      83'b?????????????????????????????????????????????????????????????????????????????1?????:
        _14951_ = b[47:40];
      83'b????????????????????????????????????????????????????????????????????????????1??????:
        _14951_ = b[55:48];
      83'b???????????????????????????????????????????????????????????????????????????1???????:
        _14951_ = b[63:56];
      83'b??????????????????????????????????????????????????????????????????????????1????????:
        _14951_ = b[71:64];
      83'b?????????????????????????????????????????????????????????????????????????1?????????:
        _14951_ = b[79:72];
      83'b????????????????????????????????????????????????????????????????????????1??????????:
        _14951_ = b[87:80];
      83'b???????????????????????????????????????????????????????????????????????1???????????:
        _14951_ = b[95:88];
      83'b??????????????????????????????????????????????????????????????????????1????????????:
        _14951_ = b[103:96];
      83'b?????????????????????????????????????????????????????????????????????1?????????????:
        _14951_ = b[111:104];
      83'b????????????????????????????????????????????????????????????????????1??????????????:
        _14951_ = b[119:112];
      83'b???????????????????????????????????????????????????????????????????1???????????????:
        _14951_ = b[127:120];
      83'b??????????????????????????????????????????????????????????????????1????????????????:
        _14951_ = b[135:128];
      83'b?????????????????????????????????????????????????????????????????1?????????????????:
        _14951_ = b[143:136];
      83'b????????????????????????????????????????????????????????????????1??????????????????:
        _14951_ = b[151:144];
      83'b???????????????????????????????????????????????????????????????1???????????????????:
        _14951_ = b[159:152];
      83'b??????????????????????????????????????????????????????????????1????????????????????:
        _14951_ = b[167:160];
      83'b?????????????????????????????????????????????????????????????1?????????????????????:
        _14951_ = b[175:168];
      83'b????????????????????????????????????????????????????????????1??????????????????????:
        _14951_ = b[183:176];
      83'b???????????????????????????????????????????????????????????1???????????????????????:
        _14951_ = b[191:184];
      83'b??????????????????????????????????????????????????????????1????????????????????????:
        _14951_ = b[199:192];
      83'b?????????????????????????????????????????????????????????1?????????????????????????:
        _14951_ = b[207:200];
      83'b????????????????????????????????????????????????????????1??????????????????????????:
        _14951_ = b[215:208];
      83'b???????????????????????????????????????????????????????1???????????????????????????:
        _14951_ = b[223:216];
      83'b??????????????????????????????????????????????????????1????????????????????????????:
        _14951_ = b[231:224];
      83'b?????????????????????????????????????????????????????1?????????????????????????????:
        _14951_ = b[239:232];
      83'b????????????????????????????????????????????????????1??????????????????????????????:
        _14951_ = b[247:240];
      83'b???????????????????????????????????????????????????1???????????????????????????????:
        _14951_ = b[255:248];
      83'b??????????????????????????????????????????????????1????????????????????????????????:
        _14951_ = b[263:256];
      83'b?????????????????????????????????????????????????1?????????????????????????????????:
        _14951_ = b[271:264];
      83'b????????????????????????????????????????????????1??????????????????????????????????:
        _14951_ = b[279:272];
      83'b???????????????????????????????????????????????1???????????????????????????????????:
        _14951_ = b[287:280];
      83'b??????????????????????????????????????????????1????????????????????????????????????:
        _14951_ = b[295:288];
      83'b?????????????????????????????????????????????1?????????????????????????????????????:
        _14951_ = b[303:296];
      83'b????????????????????????????????????????????1??????????????????????????????????????:
        _14951_ = b[311:304];
      83'b???????????????????????????????????????????1???????????????????????????????????????:
        _14951_ = b[319:312];
      83'b??????????????????????????????????????????1????????????????????????????????????????:
        _14951_ = b[327:320];
      83'b?????????????????????????????????????????1?????????????????????????????????????????:
        _14951_ = b[335:328];
      83'b????????????????????????????????????????1??????????????????????????????????????????:
        _14951_ = b[343:336];
      83'b???????????????????????????????????????1???????????????????????????????????????????:
        _14951_ = b[351:344];
      83'b??????????????????????????????????????1????????????????????????????????????????????:
        _14951_ = b[359:352];
      83'b?????????????????????????????????????1?????????????????????????????????????????????:
        _14951_ = b[367:360];
      83'b????????????????????????????????????1??????????????????????????????????????????????:
        _14951_ = b[375:368];
      83'b???????????????????????????????????1???????????????????????????????????????????????:
        _14951_ = b[383:376];
      83'b??????????????????????????????????1????????????????????????????????????????????????:
        _14951_ = b[391:384];
      83'b?????????????????????????????????1?????????????????????????????????????????????????:
        _14951_ = b[399:392];
      83'b????????????????????????????????1??????????????????????????????????????????????????:
        _14951_ = b[407:400];
      83'b???????????????????????????????1???????????????????????????????????????????????????:
        _14951_ = b[415:408];
      83'b??????????????????????????????1????????????????????????????????????????????????????:
        _14951_ = b[423:416];
      83'b?????????????????????????????1?????????????????????????????????????????????????????:
        _14951_ = b[431:424];
      83'b????????????????????????????1??????????????????????????????????????????????????????:
        _14951_ = b[439:432];
      83'b???????????????????????????1???????????????????????????????????????????????????????:
        _14951_ = b[447:440];
      83'b??????????????????????????1????????????????????????????????????????????????????????:
        _14951_ = b[455:448];
      83'b?????????????????????????1?????????????????????????????????????????????????????????:
        _14951_ = b[463:456];
      83'b????????????????????????1??????????????????????????????????????????????????????????:
        _14951_ = b[471:464];
      83'b???????????????????????1???????????????????????????????????????????????????????????:
        _14951_ = b[479:472];
      83'b??????????????????????1????????????????????????????????????????????????????????????:
        _14951_ = b[487:480];
      83'b?????????????????????1?????????????????????????????????????????????????????????????:
        _14951_ = b[495:488];
      83'b????????????????????1??????????????????????????????????????????????????????????????:
        _14951_ = b[503:496];
      83'b???????????????????1???????????????????????????????????????????????????????????????:
        _14951_ = b[511:504];
      83'b??????????????????1????????????????????????????????????????????????????????????????:
        _14951_ = b[519:512];
      83'b?????????????????1?????????????????????????????????????????????????????????????????:
        _14951_ = b[527:520];
      83'b????????????????1??????????????????????????????????????????????????????????????????:
        _14951_ = b[535:528];
      83'b???????????????1???????????????????????????????????????????????????????????????????:
        _14951_ = b[543:536];
      83'b??????????????1????????????????????????????????????????????????????????????????????:
        _14951_ = b[551:544];
      83'b?????????????1?????????????????????????????????????????????????????????????????????:
        _14951_ = b[559:552];
      83'b????????????1??????????????????????????????????????????????????????????????????????:
        _14951_ = b[567:560];
      83'b???????????1???????????????????????????????????????????????????????????????????????:
        _14951_ = b[575:568];
      83'b??????????1????????????????????????????????????????????????????????????????????????:
        _14951_ = b[583:576];
      83'b?????????1?????????????????????????????????????????????????????????????????????????:
        _14951_ = b[591:584];
      83'b????????1??????????????????????????????????????????????????????????????????????????:
        _14951_ = b[599:592];
      83'b???????1???????????????????????????????????????????????????????????????????????????:
        _14951_ = b[607:600];
      83'b??????1????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[615:608];
      83'b?????1?????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[623:616];
      83'b????1??????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[631:624];
      83'b???1???????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[639:632];
      83'b??1????????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[647:640];
      83'b?1?????????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[655:648];
      83'b1??????????????????????????????????????????????????????????????????????????????????:
        _14951_ = b[663:656];
      default:
        _14951_ = a;
    endcase
  endfunction
  assign vec_data_082 = _14951_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648], data_d1[663:656] }, { _05598_, _05597_, _05596_, _05595_, _05594_, _05593_, _05592_, _05591_, _05590_, _05589_, _05588_, _05587_, _05586_, _05585_, _05584_, _05583_, _05582_, _05581_, _05580_, _05579_, _05578_, _05577_, _05576_, _05575_, _05574_, _05573_, _05572_, _05571_, _05570_, _05569_, _05568_, _05567_, _05566_, _05565_, _05564_, _05563_, _05562_, _05561_, _05560_, _05559_, _05558_, _05557_, _05556_, _05555_, _05554_, _05553_, _05552_, _05551_, _05550_, _05549_, _05548_, _05547_, _05546_, _05545_, _05544_, _05543_, _05542_, _05541_, _05540_, _05539_, _05538_, _05537_, _05536_, _05535_, _05534_, _05533_, _05532_, _05531_, _05530_, _05529_, _05528_, _05527_, _05526_, _05525_, _05524_, _05523_, _05522_, _05521_, _05520_, _05519_, _05518_, _05517_, _05516_ });
  assign _05516_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1010011;
  assign _05517_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1010010;
  assign _05518_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1010001;
  assign _05519_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1010000;
  assign _05520_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001111;
  assign _05521_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001110;
  assign _05522_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001101;
  assign _05523_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001100;
  assign _05524_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001011;
  assign _05525_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001010;
  assign _05526_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001001;
  assign _05527_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1001000;
  assign _05528_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000111;
  assign _05529_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000110;
  assign _05530_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000101;
  assign _05531_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000100;
  assign _05532_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000011;
  assign _05533_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000010;
  assign _05534_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000001;
  assign _05535_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 7'b1000000;
  assign _05536_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111111;
  assign _05537_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111110;
  assign _05538_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111101;
  assign _05539_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111100;
  assign _05540_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111011;
  assign _05541_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111010;
  assign _05542_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111001;
  assign _05543_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b111000;
  assign _05544_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110111;
  assign _05545_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110110;
  assign _05546_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110101;
  assign _05547_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110100;
  assign _05548_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110011;
  assign _05549_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:8000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110010;
  assign _05550_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110001;
  assign _05551_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b110000;
  assign _05552_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101111;
  assign _05553_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101110;
  assign _05554_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101101;
  assign _05555_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101100;
  assign _05556_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101011;
  assign _05557_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101010;
  assign _05558_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101001;
  assign _05559_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b101000;
  assign _05560_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100111;
  assign _05561_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100110;
  assign _05562_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100101;
  assign _05563_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100100;
  assign _05564_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100011;
  assign _05565_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100010;
  assign _05566_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100001;
  assign _05567_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 6'b100000;
  assign _05568_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11111;
  assign _05569_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11110;
  assign _05570_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11101;
  assign _05571_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11100;
  assign _05572_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11011;
  assign _05573_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11010;
  assign _05574_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11001;
  assign _05575_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b11000;
  assign _05576_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10111;
  assign _05577_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10110;
  assign _05578_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10101;
  assign _05579_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10100;
  assign _05580_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10011;
  assign _05581_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10010;
  assign _05582_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10001;
  assign _05583_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 5'b10000;
  assign _05584_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1111;
  assign _05585_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1110;
  assign _05586_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1101;
  assign _05587_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1100;
  assign _05588_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1011;
  assign _05589_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1010;
  assign _05590_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1001;
  assign _05591_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 4'b1000;
  assign _05592_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 3'b111;
  assign _05593_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 3'b110;
  assign _05594_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 3'b101;
  assign _05595_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 3'b100;
  assign _05596_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 2'b11;
  assign _05597_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 2'b10;
  assign _05598_ = vec_sum_082_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7950" *) 1'b1;
  function [7:0] _15035_;
    input [7:0] a;
    input [655:0] b;
    input [81:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *)
    (* parallel_case *)
    casez (s)
      82'b?????????????????????????????????????????????????????????????????????????????????1:
        _15035_ = b[7:0];
      82'b????????????????????????????????????????????????????????????????????????????????1?:
        _15035_ = b[15:8];
      82'b???????????????????????????????????????????????????????????????????????????????1??:
        _15035_ = b[23:16];
      82'b??????????????????????????????????????????????????????????????????????????????1???:
        _15035_ = b[31:24];
      82'b?????????????????????????????????????????????????????????????????????????????1????:
        _15035_ = b[39:32];
      82'b????????????????????????????????????????????????????????????????????????????1?????:
        _15035_ = b[47:40];
      82'b???????????????????????????????????????????????????????????????????????????1??????:
        _15035_ = b[55:48];
      82'b??????????????????????????????????????????????????????????????????????????1???????:
        _15035_ = b[63:56];
      82'b?????????????????????????????????????????????????????????????????????????1????????:
        _15035_ = b[71:64];
      82'b????????????????????????????????????????????????????????????????????????1?????????:
        _15035_ = b[79:72];
      82'b???????????????????????????????????????????????????????????????????????1??????????:
        _15035_ = b[87:80];
      82'b??????????????????????????????????????????????????????????????????????1???????????:
        _15035_ = b[95:88];
      82'b?????????????????????????????????????????????????????????????????????1????????????:
        _15035_ = b[103:96];
      82'b????????????????????????????????????????????????????????????????????1?????????????:
        _15035_ = b[111:104];
      82'b???????????????????????????????????????????????????????????????????1??????????????:
        _15035_ = b[119:112];
      82'b??????????????????????????????????????????????????????????????????1???????????????:
        _15035_ = b[127:120];
      82'b?????????????????????????????????????????????????????????????????1????????????????:
        _15035_ = b[135:128];
      82'b????????????????????????????????????????????????????????????????1?????????????????:
        _15035_ = b[143:136];
      82'b???????????????????????????????????????????????????????????????1??????????????????:
        _15035_ = b[151:144];
      82'b??????????????????????????????????????????????????????????????1???????????????????:
        _15035_ = b[159:152];
      82'b?????????????????????????????????????????????????????????????1????????????????????:
        _15035_ = b[167:160];
      82'b????????????????????????????????????????????????????????????1?????????????????????:
        _15035_ = b[175:168];
      82'b???????????????????????????????????????????????????????????1??????????????????????:
        _15035_ = b[183:176];
      82'b??????????????????????????????????????????????????????????1???????????????????????:
        _15035_ = b[191:184];
      82'b?????????????????????????????????????????????????????????1????????????????????????:
        _15035_ = b[199:192];
      82'b????????????????????????????????????????????????????????1?????????????????????????:
        _15035_ = b[207:200];
      82'b???????????????????????????????????????????????????????1??????????????????????????:
        _15035_ = b[215:208];
      82'b??????????????????????????????????????????????????????1???????????????????????????:
        _15035_ = b[223:216];
      82'b?????????????????????????????????????????????????????1????????????????????????????:
        _15035_ = b[231:224];
      82'b????????????????????????????????????????????????????1?????????????????????????????:
        _15035_ = b[239:232];
      82'b???????????????????????????????????????????????????1??????????????????????????????:
        _15035_ = b[247:240];
      82'b??????????????????????????????????????????????????1???????????????????????????????:
        _15035_ = b[255:248];
      82'b?????????????????????????????????????????????????1????????????????????????????????:
        _15035_ = b[263:256];
      82'b????????????????????????????????????????????????1?????????????????????????????????:
        _15035_ = b[271:264];
      82'b???????????????????????????????????????????????1??????????????????????????????????:
        _15035_ = b[279:272];
      82'b??????????????????????????????????????????????1???????????????????????????????????:
        _15035_ = b[287:280];
      82'b?????????????????????????????????????????????1????????????????????????????????????:
        _15035_ = b[295:288];
      82'b????????????????????????????????????????????1?????????????????????????????????????:
        _15035_ = b[303:296];
      82'b???????????????????????????????????????????1??????????????????????????????????????:
        _15035_ = b[311:304];
      82'b??????????????????????????????????????????1???????????????????????????????????????:
        _15035_ = b[319:312];
      82'b?????????????????????????????????????????1????????????????????????????????????????:
        _15035_ = b[327:320];
      82'b????????????????????????????????????????1?????????????????????????????????????????:
        _15035_ = b[335:328];
      82'b???????????????????????????????????????1??????????????????????????????????????????:
        _15035_ = b[343:336];
      82'b??????????????????????????????????????1???????????????????????????????????????????:
        _15035_ = b[351:344];
      82'b?????????????????????????????????????1????????????????????????????????????????????:
        _15035_ = b[359:352];
      82'b????????????????????????????????????1?????????????????????????????????????????????:
        _15035_ = b[367:360];
      82'b???????????????????????????????????1??????????????????????????????????????????????:
        _15035_ = b[375:368];
      82'b??????????????????????????????????1???????????????????????????????????????????????:
        _15035_ = b[383:376];
      82'b?????????????????????????????????1????????????????????????????????????????????????:
        _15035_ = b[391:384];
      82'b????????????????????????????????1?????????????????????????????????????????????????:
        _15035_ = b[399:392];
      82'b???????????????????????????????1??????????????????????????????????????????????????:
        _15035_ = b[407:400];
      82'b??????????????????????????????1???????????????????????????????????????????????????:
        _15035_ = b[415:408];
      82'b?????????????????????????????1????????????????????????????????????????????????????:
        _15035_ = b[423:416];
      82'b????????????????????????????1?????????????????????????????????????????????????????:
        _15035_ = b[431:424];
      82'b???????????????????????????1??????????????????????????????????????????????????????:
        _15035_ = b[439:432];
      82'b??????????????????????????1???????????????????????????????????????????????????????:
        _15035_ = b[447:440];
      82'b?????????????????????????1????????????????????????????????????????????????????????:
        _15035_ = b[455:448];
      82'b????????????????????????1?????????????????????????????????????????????????????????:
        _15035_ = b[463:456];
      82'b???????????????????????1??????????????????????????????????????????????????????????:
        _15035_ = b[471:464];
      82'b??????????????????????1???????????????????????????????????????????????????????????:
        _15035_ = b[479:472];
      82'b?????????????????????1????????????????????????????????????????????????????????????:
        _15035_ = b[487:480];
      82'b????????????????????1?????????????????????????????????????????????????????????????:
        _15035_ = b[495:488];
      82'b???????????????????1??????????????????????????????????????????????????????????????:
        _15035_ = b[503:496];
      82'b??????????????????1???????????????????????????????????????????????????????????????:
        _15035_ = b[511:504];
      82'b?????????????????1????????????????????????????????????????????????????????????????:
        _15035_ = b[519:512];
      82'b????????????????1?????????????????????????????????????????????????????????????????:
        _15035_ = b[527:520];
      82'b???????????????1??????????????????????????????????????????????????????????????????:
        _15035_ = b[535:528];
      82'b??????????????1???????????????????????????????????????????????????????????????????:
        _15035_ = b[543:536];
      82'b?????????????1????????????????????????????????????????????????????????????????????:
        _15035_ = b[551:544];
      82'b????????????1?????????????????????????????????????????????????????????????????????:
        _15035_ = b[559:552];
      82'b???????????1??????????????????????????????????????????????????????????????????????:
        _15035_ = b[567:560];
      82'b??????????1???????????????????????????????????????????????????????????????????????:
        _15035_ = b[575:568];
      82'b?????????1????????????????????????????????????????????????????????????????????????:
        _15035_ = b[583:576];
      82'b????????1?????????????????????????????????????????????????????????????????????????:
        _15035_ = b[591:584];
      82'b???????1??????????????????????????????????????????????????????????????????????????:
        _15035_ = b[599:592];
      82'b??????1???????????????????????????????????????????????????????????????????????????:
        _15035_ = b[607:600];
      82'b?????1????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[615:608];
      82'b????1?????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[623:616];
      82'b???1??????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[631:624];
      82'b??1???????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[639:632];
      82'b?1????????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[647:640];
      82'b1?????????????????????????????????????????????????????????????????????????????????:
        _15035_ = b[655:648];
      default:
        _15035_ = a;
    endcase
  endfunction
  assign vec_data_081 = _15035_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640], data_d1[655:648] }, { _05680_, _05679_, _05678_, _05677_, _05676_, _05675_, _05674_, _05673_, _05672_, _05671_, _05670_, _05669_, _05668_, _05667_, _05666_, _05665_, _05664_, _05663_, _05662_, _05661_, _05660_, _05659_, _05658_, _05657_, _05656_, _05655_, _05654_, _05653_, _05652_, _05651_, _05650_, _05649_, _05648_, _05647_, _05646_, _05645_, _05644_, _05643_, _05642_, _05641_, _05640_, _05639_, _05638_, _05637_, _05636_, _05635_, _05634_, _05633_, _05632_, _05631_, _05630_, _05629_, _05628_, _05627_, _05626_, _05625_, _05624_, _05623_, _05622_, _05621_, _05620_, _05619_, _05618_, _05617_, _05616_, _05615_, _05614_, _05613_, _05612_, _05611_, _05610_, _05609_, _05608_, _05607_, _05606_, _05605_, _05604_, _05603_, _05602_, _05601_, _05600_, _05599_ });
  assign _05599_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1010010;
  assign _05600_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1010001;
  assign _05601_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1010000;
  assign _05602_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001111;
  assign _05603_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001110;
  assign _05604_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001101;
  assign _05605_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001100;
  assign _05606_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001011;
  assign _05607_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001010;
  assign _05608_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7933|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001001;
  assign _05609_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7932|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1001000;
  assign _05610_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7931|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000111;
  assign _05611_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7930|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000110;
  assign _05612_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7929|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000101;
  assign _05613_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000100;
  assign _05614_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000011;
  assign _05615_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000010;
  assign _05616_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000001;
  assign _05617_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 7'b1000000;
  assign _05618_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111111;
  assign _05619_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111110;
  assign _05620_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111101;
  assign _05621_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111100;
  assign _05622_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111011;
  assign _05623_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111010;
  assign _05624_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111001;
  assign _05625_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b111000;
  assign _05626_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110111;
  assign _05627_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110110;
  assign _05628_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110101;
  assign _05629_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110100;
  assign _05630_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110011;
  assign _05631_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110010;
  assign _05632_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110001;
  assign _05633_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b110000;
  assign _05634_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101111;
  assign _05635_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101110;
  assign _05636_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101101;
  assign _05637_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101100;
  assign _05638_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101011;
  assign _05639_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101010;
  assign _05640_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101001;
  assign _05641_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b101000;
  assign _05642_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100111;
  assign _05643_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100110;
  assign _05644_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100101;
  assign _05645_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100100;
  assign _05646_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100011;
  assign _05647_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100010;
  assign _05648_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100001;
  assign _05649_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 6'b100000;
  assign _05650_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11111;
  assign _05651_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11110;
  assign _05652_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11101;
  assign _05653_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11100;
  assign _05654_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11011;
  assign _05655_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11010;
  assign _05656_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11001;
  assign _05657_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b11000;
  assign _05658_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10111;
  assign _05659_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10110;
  assign _05660_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10101;
  assign _05661_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10100;
  assign _05662_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10011;
  assign _05663_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10010;
  assign _05664_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10001;
  assign _05665_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 5'b10000;
  assign _05666_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1111;
  assign _05667_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1110;
  assign _05668_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1101;
  assign _05669_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1100;
  assign _05670_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1011;
  assign _05671_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1010;
  assign _05672_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1001;
  assign _05673_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 4'b1000;
  assign _05674_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 3'b111;
  assign _05675_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 3'b110;
  assign _05676_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 3'b101;
  assign _05677_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 3'b100;
  assign _05678_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 2'b11;
  assign _05679_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 2'b10;
  assign _05680_ = vec_sum_081_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7860" *) 1'b1;
  function [7:0] _15118_;
    input [7:0] a;
    input [647:0] b;
    input [80:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *)
    (* parallel_case *)
    casez (s)
      81'b????????????????????????????????????????????????????????????????????????????????1:
        _15118_ = b[7:0];
      81'b???????????????????????????????????????????????????????????????????????????????1?:
        _15118_ = b[15:8];
      81'b??????????????????????????????????????????????????????????????????????????????1??:
        _15118_ = b[23:16];
      81'b?????????????????????????????????????????????????????????????????????????????1???:
        _15118_ = b[31:24];
      81'b????????????????????????????????????????????????????????????????????????????1????:
        _15118_ = b[39:32];
      81'b???????????????????????????????????????????????????????????????????????????1?????:
        _15118_ = b[47:40];
      81'b??????????????????????????????????????????????????????????????????????????1??????:
        _15118_ = b[55:48];
      81'b?????????????????????????????????????????????????????????????????????????1???????:
        _15118_ = b[63:56];
      81'b????????????????????????????????????????????????????????????????????????1????????:
        _15118_ = b[71:64];
      81'b???????????????????????????????????????????????????????????????????????1?????????:
        _15118_ = b[79:72];
      81'b??????????????????????????????????????????????????????????????????????1??????????:
        _15118_ = b[87:80];
      81'b?????????????????????????????????????????????????????????????????????1???????????:
        _15118_ = b[95:88];
      81'b????????????????????????????????????????????????????????????????????1????????????:
        _15118_ = b[103:96];
      81'b???????????????????????????????????????????????????????????????????1?????????????:
        _15118_ = b[111:104];
      81'b??????????????????????????????????????????????????????????????????1??????????????:
        _15118_ = b[119:112];
      81'b?????????????????????????????????????????????????????????????????1???????????????:
        _15118_ = b[127:120];
      81'b????????????????????????????????????????????????????????????????1????????????????:
        _15118_ = b[135:128];
      81'b???????????????????????????????????????????????????????????????1?????????????????:
        _15118_ = b[143:136];
      81'b??????????????????????????????????????????????????????????????1??????????????????:
        _15118_ = b[151:144];
      81'b?????????????????????????????????????????????????????????????1???????????????????:
        _15118_ = b[159:152];
      81'b????????????????????????????????????????????????????????????1????????????????????:
        _15118_ = b[167:160];
      81'b???????????????????????????????????????????????????????????1?????????????????????:
        _15118_ = b[175:168];
      81'b??????????????????????????????????????????????????????????1??????????????????????:
        _15118_ = b[183:176];
      81'b?????????????????????????????????????????????????????????1???????????????????????:
        _15118_ = b[191:184];
      81'b????????????????????????????????????????????????????????1????????????????????????:
        _15118_ = b[199:192];
      81'b???????????????????????????????????????????????????????1?????????????????????????:
        _15118_ = b[207:200];
      81'b??????????????????????????????????????????????????????1??????????????????????????:
        _15118_ = b[215:208];
      81'b?????????????????????????????????????????????????????1???????????????????????????:
        _15118_ = b[223:216];
      81'b????????????????????????????????????????????????????1????????????????????????????:
        _15118_ = b[231:224];
      81'b???????????????????????????????????????????????????1?????????????????????????????:
        _15118_ = b[239:232];
      81'b??????????????????????????????????????????????????1??????????????????????????????:
        _15118_ = b[247:240];
      81'b?????????????????????????????????????????????????1???????????????????????????????:
        _15118_ = b[255:248];
      81'b????????????????????????????????????????????????1????????????????????????????????:
        _15118_ = b[263:256];
      81'b???????????????????????????????????????????????1?????????????????????????????????:
        _15118_ = b[271:264];
      81'b??????????????????????????????????????????????1??????????????????????????????????:
        _15118_ = b[279:272];
      81'b?????????????????????????????????????????????1???????????????????????????????????:
        _15118_ = b[287:280];
      81'b????????????????????????????????????????????1????????????????????????????????????:
        _15118_ = b[295:288];
      81'b???????????????????????????????????????????1?????????????????????????????????????:
        _15118_ = b[303:296];
      81'b??????????????????????????????????????????1??????????????????????????????????????:
        _15118_ = b[311:304];
      81'b?????????????????????????????????????????1???????????????????????????????????????:
        _15118_ = b[319:312];
      81'b????????????????????????????????????????1????????????????????????????????????????:
        _15118_ = b[327:320];
      81'b???????????????????????????????????????1?????????????????????????????????????????:
        _15118_ = b[335:328];
      81'b??????????????????????????????????????1??????????????????????????????????????????:
        _15118_ = b[343:336];
      81'b?????????????????????????????????????1???????????????????????????????????????????:
        _15118_ = b[351:344];
      81'b????????????????????????????????????1????????????????????????????????????????????:
        _15118_ = b[359:352];
      81'b???????????????????????????????????1?????????????????????????????????????????????:
        _15118_ = b[367:360];
      81'b??????????????????????????????????1??????????????????????????????????????????????:
        _15118_ = b[375:368];
      81'b?????????????????????????????????1???????????????????????????????????????????????:
        _15118_ = b[383:376];
      81'b????????????????????????????????1????????????????????????????????????????????????:
        _15118_ = b[391:384];
      81'b???????????????????????????????1?????????????????????????????????????????????????:
        _15118_ = b[399:392];
      81'b??????????????????????????????1??????????????????????????????????????????????????:
        _15118_ = b[407:400];
      81'b?????????????????????????????1???????????????????????????????????????????????????:
        _15118_ = b[415:408];
      81'b????????????????????????????1????????????????????????????????????????????????????:
        _15118_ = b[423:416];
      81'b???????????????????????????1?????????????????????????????????????????????????????:
        _15118_ = b[431:424];
      81'b??????????????????????????1??????????????????????????????????????????????????????:
        _15118_ = b[439:432];
      81'b?????????????????????????1???????????????????????????????????????????????????????:
        _15118_ = b[447:440];
      81'b????????????????????????1????????????????????????????????????????????????????????:
        _15118_ = b[455:448];
      81'b???????????????????????1?????????????????????????????????????????????????????????:
        _15118_ = b[463:456];
      81'b??????????????????????1??????????????????????????????????????????????????????????:
        _15118_ = b[471:464];
      81'b?????????????????????1???????????????????????????????????????????????????????????:
        _15118_ = b[479:472];
      81'b????????????????????1????????????????????????????????????????????????????????????:
        _15118_ = b[487:480];
      81'b???????????????????1?????????????????????????????????????????????????????????????:
        _15118_ = b[495:488];
      81'b??????????????????1??????????????????????????????????????????????????????????????:
        _15118_ = b[503:496];
      81'b?????????????????1???????????????????????????????????????????????????????????????:
        _15118_ = b[511:504];
      81'b????????????????1????????????????????????????????????????????????????????????????:
        _15118_ = b[519:512];
      81'b???????????????1?????????????????????????????????????????????????????????????????:
        _15118_ = b[527:520];
      81'b??????????????1??????????????????????????????????????????????????????????????????:
        _15118_ = b[535:528];
      81'b?????????????1???????????????????????????????????????????????????????????????????:
        _15118_ = b[543:536];
      81'b????????????1????????????????????????????????????????????????????????????????????:
        _15118_ = b[551:544];
      81'b???????????1?????????????????????????????????????????????????????????????????????:
        _15118_ = b[559:552];
      81'b??????????1??????????????????????????????????????????????????????????????????????:
        _15118_ = b[567:560];
      81'b?????????1???????????????????????????????????????????????????????????????????????:
        _15118_ = b[575:568];
      81'b????????1????????????????????????????????????????????????????????????????????????:
        _15118_ = b[583:576];
      81'b???????1?????????????????????????????????????????????????????????????????????????:
        _15118_ = b[591:584];
      81'b??????1??????????????????????????????????????????????????????????????????????????:
        _15118_ = b[599:592];
      81'b?????1???????????????????????????????????????????????????????????????????????????:
        _15118_ = b[607:600];
      81'b????1????????????????????????????????????????????????????????????????????????????:
        _15118_ = b[615:608];
      81'b???1?????????????????????????????????????????????????????????????????????????????:
        _15118_ = b[623:616];
      81'b??1??????????????????????????????????????????????????????????????????????????????:
        _15118_ = b[631:624];
      81'b?1???????????????????????????????????????????????????????????????????????????????:
        _15118_ = b[639:632];
      81'b1????????????????????????????????????????????????????????????????????????????????:
        _15118_ = b[647:640];
      default:
        _15118_ = a;
    endcase
  endfunction
  assign vec_data_080 = _15118_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632], data_d1[647:640] }, { _05761_, _05760_, _05759_, _05758_, _05757_, _05756_, _05755_, _05754_, _05753_, _05752_, _05751_, _05750_, _05749_, _05748_, _05747_, _05746_, _05745_, _05744_, _05743_, _05742_, _05741_, _05740_, _05739_, _05738_, _05737_, _05736_, _05735_, _05734_, _05733_, _05732_, _05731_, _05730_, _05729_, _05728_, _05727_, _05726_, _05725_, _05724_, _05723_, _05722_, _05721_, _05720_, _05719_, _05718_, _05717_, _05716_, _05715_, _05714_, _05713_, _05712_, _05711_, _05710_, _05709_, _05708_, _05707_, _05706_, _05705_, _05704_, _05703_, _05702_, _05701_, _05700_, _05699_, _05698_, _05697_, _05696_, _05695_, _05694_, _05693_, _05692_, _05691_, _05690_, _05689_, _05688_, _05687_, _05686_, _05685_, _05684_, _05683_, _05682_, _05681_ });
  assign _05681_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1010001;
  assign _05682_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1010000;
  assign _05683_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001111;
  assign _05684_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001110;
  assign _05685_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001101;
  assign _05686_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001100;
  assign _05687_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001011;
  assign _05688_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001010;
  assign _05689_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001001;
  assign _05690_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1001000;
  assign _05691_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000111;
  assign _05692_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000110;
  assign _05693_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000101;
  assign _05694_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000100;
  assign _05695_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000011;
  assign _05696_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000010;
  assign _05697_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000001;
  assign _05698_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 7'b1000000;
  assign _05699_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111111;
  assign _05700_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111110;
  assign _05701_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111101;
  assign _05702_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111100;
  assign _05703_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111011;
  assign _05704_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111010;
  assign _05705_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111001;
  assign _05706_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b111000;
  assign _05707_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110111;
  assign _05708_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110110;
  assign _05709_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110101;
  assign _05710_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110100;
  assign _05711_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110011;
  assign _05712_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110010;
  assign _05713_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110001;
  assign _05714_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b110000;
  assign _05715_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101111;
  assign _05716_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101110;
  assign _05717_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101101;
  assign _05718_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101100;
  assign _05719_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101011;
  assign _05720_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101010;
  assign _05721_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101001;
  assign _05722_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b101000;
  assign _05723_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100111;
  assign _05724_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100110;
  assign _05725_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100101;
  assign _05726_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100100;
  assign _05727_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100011;
  assign _05728_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100010;
  assign _05729_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100001;
  assign _05730_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 6'b100000;
  assign _05731_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11111;
  assign _05732_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11110;
  assign _05733_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11101;
  assign _05734_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11100;
  assign _05735_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11011;
  assign _05736_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11010;
  assign _05737_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11001;
  assign _05738_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b11000;
  assign _05739_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10111;
  assign _05740_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10110;
  assign _05741_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10101;
  assign _05742_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10100;
  assign _05743_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10011;
  assign _05744_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10010;
  assign _05745_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10001;
  assign _05746_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 5'b10000;
  assign _05747_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1111;
  assign _05748_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1110;
  assign _05749_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1101;
  assign _05750_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1100;
  assign _05751_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1011;
  assign _05752_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1010;
  assign _05753_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1001;
  assign _05754_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 4'b1000;
  assign _05755_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 3'b111;
  assign _05756_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 3'b110;
  assign _05757_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 3'b101;
  assign _05758_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 3'b100;
  assign _05759_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 2'b11;
  assign _05760_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 2'b10;
  assign _05761_ = vec_sum_080_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7771" *) 1'b1;
  function [7:0] _15200_;
    input [7:0] a;
    input [639:0] b;
    input [79:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *)
    (* parallel_case *)
    casez (s)
      80'b???????????????????????????????????????????????????????????????????????????????1:
        _15200_ = b[7:0];
      80'b??????????????????????????????????????????????????????????????????????????????1?:
        _15200_ = b[15:8];
      80'b?????????????????????????????????????????????????????????????????????????????1??:
        _15200_ = b[23:16];
      80'b????????????????????????????????????????????????????????????????????????????1???:
        _15200_ = b[31:24];
      80'b???????????????????????????????????????????????????????????????????????????1????:
        _15200_ = b[39:32];
      80'b??????????????????????????????????????????????????????????????????????????1?????:
        _15200_ = b[47:40];
      80'b?????????????????????????????????????????????????????????????????????????1??????:
        _15200_ = b[55:48];
      80'b????????????????????????????????????????????????????????????????????????1???????:
        _15200_ = b[63:56];
      80'b???????????????????????????????????????????????????????????????????????1????????:
        _15200_ = b[71:64];
      80'b??????????????????????????????????????????????????????????????????????1?????????:
        _15200_ = b[79:72];
      80'b?????????????????????????????????????????????????????????????????????1??????????:
        _15200_ = b[87:80];
      80'b????????????????????????????????????????????????????????????????????1???????????:
        _15200_ = b[95:88];
      80'b???????????????????????????????????????????????????????????????????1????????????:
        _15200_ = b[103:96];
      80'b??????????????????????????????????????????????????????????????????1?????????????:
        _15200_ = b[111:104];
      80'b?????????????????????????????????????????????????????????????????1??????????????:
        _15200_ = b[119:112];
      80'b????????????????????????????????????????????????????????????????1???????????????:
        _15200_ = b[127:120];
      80'b???????????????????????????????????????????????????????????????1????????????????:
        _15200_ = b[135:128];
      80'b??????????????????????????????????????????????????????????????1?????????????????:
        _15200_ = b[143:136];
      80'b?????????????????????????????????????????????????????????????1??????????????????:
        _15200_ = b[151:144];
      80'b????????????????????????????????????????????????????????????1???????????????????:
        _15200_ = b[159:152];
      80'b???????????????????????????????????????????????????????????1????????????????????:
        _15200_ = b[167:160];
      80'b??????????????????????????????????????????????????????????1?????????????????????:
        _15200_ = b[175:168];
      80'b?????????????????????????????????????????????????????????1??????????????????????:
        _15200_ = b[183:176];
      80'b????????????????????????????????????????????????????????1???????????????????????:
        _15200_ = b[191:184];
      80'b???????????????????????????????????????????????????????1????????????????????????:
        _15200_ = b[199:192];
      80'b??????????????????????????????????????????????????????1?????????????????????????:
        _15200_ = b[207:200];
      80'b?????????????????????????????????????????????????????1??????????????????????????:
        _15200_ = b[215:208];
      80'b????????????????????????????????????????????????????1???????????????????????????:
        _15200_ = b[223:216];
      80'b???????????????????????????????????????????????????1????????????????????????????:
        _15200_ = b[231:224];
      80'b??????????????????????????????????????????????????1?????????????????????????????:
        _15200_ = b[239:232];
      80'b?????????????????????????????????????????????????1??????????????????????????????:
        _15200_ = b[247:240];
      80'b????????????????????????????????????????????????1???????????????????????????????:
        _15200_ = b[255:248];
      80'b???????????????????????????????????????????????1????????????????????????????????:
        _15200_ = b[263:256];
      80'b??????????????????????????????????????????????1?????????????????????????????????:
        _15200_ = b[271:264];
      80'b?????????????????????????????????????????????1??????????????????????????????????:
        _15200_ = b[279:272];
      80'b????????????????????????????????????????????1???????????????????????????????????:
        _15200_ = b[287:280];
      80'b???????????????????????????????????????????1????????????????????????????????????:
        _15200_ = b[295:288];
      80'b??????????????????????????????????????????1?????????????????????????????????????:
        _15200_ = b[303:296];
      80'b?????????????????????????????????????????1??????????????????????????????????????:
        _15200_ = b[311:304];
      80'b????????????????????????????????????????1???????????????????????????????????????:
        _15200_ = b[319:312];
      80'b???????????????????????????????????????1????????????????????????????????????????:
        _15200_ = b[327:320];
      80'b??????????????????????????????????????1?????????????????????????????????????????:
        _15200_ = b[335:328];
      80'b?????????????????????????????????????1??????????????????????????????????????????:
        _15200_ = b[343:336];
      80'b????????????????????????????????????1???????????????????????????????????????????:
        _15200_ = b[351:344];
      80'b???????????????????????????????????1????????????????????????????????????????????:
        _15200_ = b[359:352];
      80'b??????????????????????????????????1?????????????????????????????????????????????:
        _15200_ = b[367:360];
      80'b?????????????????????????????????1??????????????????????????????????????????????:
        _15200_ = b[375:368];
      80'b????????????????????????????????1???????????????????????????????????????????????:
        _15200_ = b[383:376];
      80'b???????????????????????????????1????????????????????????????????????????????????:
        _15200_ = b[391:384];
      80'b??????????????????????????????1?????????????????????????????????????????????????:
        _15200_ = b[399:392];
      80'b?????????????????????????????1??????????????????????????????????????????????????:
        _15200_ = b[407:400];
      80'b????????????????????????????1???????????????????????????????????????????????????:
        _15200_ = b[415:408];
      80'b???????????????????????????1????????????????????????????????????????????????????:
        _15200_ = b[423:416];
      80'b??????????????????????????1?????????????????????????????????????????????????????:
        _15200_ = b[431:424];
      80'b?????????????????????????1??????????????????????????????????????????????????????:
        _15200_ = b[439:432];
      80'b????????????????????????1???????????????????????????????????????????????????????:
        _15200_ = b[447:440];
      80'b???????????????????????1????????????????????????????????????????????????????????:
        _15200_ = b[455:448];
      80'b??????????????????????1?????????????????????????????????????????????????????????:
        _15200_ = b[463:456];
      80'b?????????????????????1??????????????????????????????????????????????????????????:
        _15200_ = b[471:464];
      80'b????????????????????1???????????????????????????????????????????????????????????:
        _15200_ = b[479:472];
      80'b???????????????????1????????????????????????????????????????????????????????????:
        _15200_ = b[487:480];
      80'b??????????????????1?????????????????????????????????????????????????????????????:
        _15200_ = b[495:488];
      80'b?????????????????1??????????????????????????????????????????????????????????????:
        _15200_ = b[503:496];
      80'b????????????????1???????????????????????????????????????????????????????????????:
        _15200_ = b[511:504];
      80'b???????????????1????????????????????????????????????????????????????????????????:
        _15200_ = b[519:512];
      80'b??????????????1?????????????????????????????????????????????????????????????????:
        _15200_ = b[527:520];
      80'b?????????????1??????????????????????????????????????????????????????????????????:
        _15200_ = b[535:528];
      80'b????????????1???????????????????????????????????????????????????????????????????:
        _15200_ = b[543:536];
      80'b???????????1????????????????????????????????????????????????????????????????????:
        _15200_ = b[551:544];
      80'b??????????1?????????????????????????????????????????????????????????????????????:
        _15200_ = b[559:552];
      80'b?????????1??????????????????????????????????????????????????????????????????????:
        _15200_ = b[567:560];
      80'b????????1???????????????????????????????????????????????????????????????????????:
        _15200_ = b[575:568];
      80'b???????1????????????????????????????????????????????????????????????????????????:
        _15200_ = b[583:576];
      80'b??????1?????????????????????????????????????????????????????????????????????????:
        _15200_ = b[591:584];
      80'b?????1??????????????????????????????????????????????????????????????????????????:
        _15200_ = b[599:592];
      80'b????1???????????????????????????????????????????????????????????????????????????:
        _15200_ = b[607:600];
      80'b???1????????????????????????????????????????????????????????????????????????????:
        _15200_ = b[615:608];
      80'b??1?????????????????????????????????????????????????????????????????????????????:
        _15200_ = b[623:616];
      80'b?1??????????????????????????????????????????????????????????????????????????????:
        _15200_ = b[631:624];
      80'b1???????????????????????????????????????????????????????????????????????????????:
        _15200_ = b[639:632];
      default:
        _15200_ = a;
    endcase
  endfunction
  assign vec_data_079 = _15200_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624], data_d1[639:632] }, { _05841_, _05840_, _05839_, _05838_, _05837_, _05836_, _05835_, _05834_, _05833_, _05832_, _05831_, _05830_, _05829_, _05828_, _05827_, _05826_, _05825_, _05824_, _05823_, _05822_, _05821_, _05820_, _05819_, _05818_, _05817_, _05816_, _05815_, _05814_, _05813_, _05812_, _05811_, _05810_, _05809_, _05808_, _05807_, _05806_, _05805_, _05804_, _05803_, _05802_, _05801_, _05800_, _05799_, _05798_, _05797_, _05796_, _05795_, _05794_, _05793_, _05792_, _05791_, _05790_, _05789_, _05788_, _05787_, _05786_, _05785_, _05784_, _05783_, _05782_, _05781_, _05780_, _05779_, _05778_, _05777_, _05776_, _05775_, _05774_, _05773_, _05772_, _05771_, _05770_, _05769_, _05768_, _05767_, _05766_, _05765_, _05764_, _05763_, _05762_ });
  assign _05762_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1010000;
  assign _05763_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001111;
  assign _05764_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001110;
  assign _05765_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001101;
  assign _05766_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001100;
  assign _05767_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001011;
  assign _05768_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001010;
  assign _05769_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001001;
  assign _05770_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1001000;
  assign _05771_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000111;
  assign _05772_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000110;
  assign _05773_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000101;
  assign _05774_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000100;
  assign _05775_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000011;
  assign _05776_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000010;
  assign _05777_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000001;
  assign _05778_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 7'b1000000;
  assign _05779_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111111;
  assign _05780_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111110;
  assign _05781_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111101;
  assign _05782_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111100;
  assign _05783_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111011;
  assign _05784_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111010;
  assign _05785_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111001;
  assign _05786_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b111000;
  assign _05787_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110111;
  assign _05788_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110110;
  assign _05789_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110101;
  assign _05790_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110100;
  assign _05791_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110011;
  assign _05792_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110010;
  assign _05793_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110001;
  assign _05794_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b110000;
  assign _05795_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101111;
  assign _05796_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101110;
  assign _05797_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101101;
  assign _05798_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101100;
  assign _05799_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101011;
  assign _05800_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101010;
  assign _05801_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101001;
  assign _05802_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b101000;
  assign _05803_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100111;
  assign _05804_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100110;
  assign _05805_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100101;
  assign _05806_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100100;
  assign _05807_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100011;
  assign _05808_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100010;
  assign _05809_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100001;
  assign _05810_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 6'b100000;
  assign _05811_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11111;
  assign _05812_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11110;
  assign _05813_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11101;
  assign _05814_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11100;
  assign _05815_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11011;
  assign _05816_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11010;
  assign _05817_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11001;
  assign _05818_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b11000;
  assign _05819_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10111;
  assign _05820_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10110;
  assign _05821_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10101;
  assign _05822_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10100;
  assign _05823_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10011;
  assign _05824_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10010;
  assign _05825_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10001;
  assign _05826_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 5'b10000;
  assign _05827_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1111;
  assign _05828_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1110;
  assign _05829_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1101;
  assign _05830_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1100;
  assign _05831_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1011;
  assign _05832_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1010;
  assign _05833_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1001;
  assign _05834_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 4'b1000;
  assign _05835_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 3'b111;
  assign _05836_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 3'b110;
  assign _05837_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 3'b101;
  assign _05838_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 3'b100;
  assign _05839_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 2'b11;
  assign _05840_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 2'b10;
  assign _05841_ = vec_sum_079_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7683" *) 1'b1;
  function [7:0] _15281_;
    input [7:0] a;
    input [631:0] b;
    input [78:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *)
    (* parallel_case *)
    casez (s)
      79'b??????????????????????????????????????????????????????????????????????????????1:
        _15281_ = b[7:0];
      79'b?????????????????????????????????????????????????????????????????????????????1?:
        _15281_ = b[15:8];
      79'b????????????????????????????????????????????????????????????????????????????1??:
        _15281_ = b[23:16];
      79'b???????????????????????????????????????????????????????????????????????????1???:
        _15281_ = b[31:24];
      79'b??????????????????????????????????????????????????????????????????????????1????:
        _15281_ = b[39:32];
      79'b?????????????????????????????????????????????????????????????????????????1?????:
        _15281_ = b[47:40];
      79'b????????????????????????????????????????????????????????????????????????1??????:
        _15281_ = b[55:48];
      79'b???????????????????????????????????????????????????????????????????????1???????:
        _15281_ = b[63:56];
      79'b??????????????????????????????????????????????????????????????????????1????????:
        _15281_ = b[71:64];
      79'b?????????????????????????????????????????????????????????????????????1?????????:
        _15281_ = b[79:72];
      79'b????????????????????????????????????????????????????????????????????1??????????:
        _15281_ = b[87:80];
      79'b???????????????????????????????????????????????????????????????????1???????????:
        _15281_ = b[95:88];
      79'b??????????????????????????????????????????????????????????????????1????????????:
        _15281_ = b[103:96];
      79'b?????????????????????????????????????????????????????????????????1?????????????:
        _15281_ = b[111:104];
      79'b????????????????????????????????????????????????????????????????1??????????????:
        _15281_ = b[119:112];
      79'b???????????????????????????????????????????????????????????????1???????????????:
        _15281_ = b[127:120];
      79'b??????????????????????????????????????????????????????????????1????????????????:
        _15281_ = b[135:128];
      79'b?????????????????????????????????????????????????????????????1?????????????????:
        _15281_ = b[143:136];
      79'b????????????????????????????????????????????????????????????1??????????????????:
        _15281_ = b[151:144];
      79'b???????????????????????????????????????????????????????????1???????????????????:
        _15281_ = b[159:152];
      79'b??????????????????????????????????????????????????????????1????????????????????:
        _15281_ = b[167:160];
      79'b?????????????????????????????????????????????????????????1?????????????????????:
        _15281_ = b[175:168];
      79'b????????????????????????????????????????????????????????1??????????????????????:
        _15281_ = b[183:176];
      79'b???????????????????????????????????????????????????????1???????????????????????:
        _15281_ = b[191:184];
      79'b??????????????????????????????????????????????????????1????????????????????????:
        _15281_ = b[199:192];
      79'b?????????????????????????????????????????????????????1?????????????????????????:
        _15281_ = b[207:200];
      79'b????????????????????????????????????????????????????1??????????????????????????:
        _15281_ = b[215:208];
      79'b???????????????????????????????????????????????????1???????????????????????????:
        _15281_ = b[223:216];
      79'b??????????????????????????????????????????????????1????????????????????????????:
        _15281_ = b[231:224];
      79'b?????????????????????????????????????????????????1?????????????????????????????:
        _15281_ = b[239:232];
      79'b????????????????????????????????????????????????1??????????????????????????????:
        _15281_ = b[247:240];
      79'b???????????????????????????????????????????????1???????????????????????????????:
        _15281_ = b[255:248];
      79'b??????????????????????????????????????????????1????????????????????????????????:
        _15281_ = b[263:256];
      79'b?????????????????????????????????????????????1?????????????????????????????????:
        _15281_ = b[271:264];
      79'b????????????????????????????????????????????1??????????????????????????????????:
        _15281_ = b[279:272];
      79'b???????????????????????????????????????????1???????????????????????????????????:
        _15281_ = b[287:280];
      79'b??????????????????????????????????????????1????????????????????????????????????:
        _15281_ = b[295:288];
      79'b?????????????????????????????????????????1?????????????????????????????????????:
        _15281_ = b[303:296];
      79'b????????????????????????????????????????1??????????????????????????????????????:
        _15281_ = b[311:304];
      79'b???????????????????????????????????????1???????????????????????????????????????:
        _15281_ = b[319:312];
      79'b??????????????????????????????????????1????????????????????????????????????????:
        _15281_ = b[327:320];
      79'b?????????????????????????????????????1?????????????????????????????????????????:
        _15281_ = b[335:328];
      79'b????????????????????????????????????1??????????????????????????????????????????:
        _15281_ = b[343:336];
      79'b???????????????????????????????????1???????????????????????????????????????????:
        _15281_ = b[351:344];
      79'b??????????????????????????????????1????????????????????????????????????????????:
        _15281_ = b[359:352];
      79'b?????????????????????????????????1?????????????????????????????????????????????:
        _15281_ = b[367:360];
      79'b????????????????????????????????1??????????????????????????????????????????????:
        _15281_ = b[375:368];
      79'b???????????????????????????????1???????????????????????????????????????????????:
        _15281_ = b[383:376];
      79'b??????????????????????????????1????????????????????????????????????????????????:
        _15281_ = b[391:384];
      79'b?????????????????????????????1?????????????????????????????????????????????????:
        _15281_ = b[399:392];
      79'b????????????????????????????1??????????????????????????????????????????????????:
        _15281_ = b[407:400];
      79'b???????????????????????????1???????????????????????????????????????????????????:
        _15281_ = b[415:408];
      79'b??????????????????????????1????????????????????????????????????????????????????:
        _15281_ = b[423:416];
      79'b?????????????????????????1?????????????????????????????????????????????????????:
        _15281_ = b[431:424];
      79'b????????????????????????1??????????????????????????????????????????????????????:
        _15281_ = b[439:432];
      79'b???????????????????????1???????????????????????????????????????????????????????:
        _15281_ = b[447:440];
      79'b??????????????????????1????????????????????????????????????????????????????????:
        _15281_ = b[455:448];
      79'b?????????????????????1?????????????????????????????????????????????????????????:
        _15281_ = b[463:456];
      79'b????????????????????1??????????????????????????????????????????????????????????:
        _15281_ = b[471:464];
      79'b???????????????????1???????????????????????????????????????????????????????????:
        _15281_ = b[479:472];
      79'b??????????????????1????????????????????????????????????????????????????????????:
        _15281_ = b[487:480];
      79'b?????????????????1?????????????????????????????????????????????????????????????:
        _15281_ = b[495:488];
      79'b????????????????1??????????????????????????????????????????????????????????????:
        _15281_ = b[503:496];
      79'b???????????????1???????????????????????????????????????????????????????????????:
        _15281_ = b[511:504];
      79'b??????????????1????????????????????????????????????????????????????????????????:
        _15281_ = b[519:512];
      79'b?????????????1?????????????????????????????????????????????????????????????????:
        _15281_ = b[527:520];
      79'b????????????1??????????????????????????????????????????????????????????????????:
        _15281_ = b[535:528];
      79'b???????????1???????????????????????????????????????????????????????????????????:
        _15281_ = b[543:536];
      79'b??????????1????????????????????????????????????????????????????????????????????:
        _15281_ = b[551:544];
      79'b?????????1?????????????????????????????????????????????????????????????????????:
        _15281_ = b[559:552];
      79'b????????1??????????????????????????????????????????????????????????????????????:
        _15281_ = b[567:560];
      79'b???????1???????????????????????????????????????????????????????????????????????:
        _15281_ = b[575:568];
      79'b??????1????????????????????????????????????????????????????????????????????????:
        _15281_ = b[583:576];
      79'b?????1?????????????????????????????????????????????????????????????????????????:
        _15281_ = b[591:584];
      79'b????1??????????????????????????????????????????????????????????????????????????:
        _15281_ = b[599:592];
      79'b???1???????????????????????????????????????????????????????????????????????????:
        _15281_ = b[607:600];
      79'b??1????????????????????????????????????????????????????????????????????????????:
        _15281_ = b[615:608];
      79'b?1?????????????????????????????????????????????????????????????????????????????:
        _15281_ = b[623:616];
      79'b1??????????????????????????????????????????????????????????????????????????????:
        _15281_ = b[631:624];
      default:
        _15281_ = a;
    endcase
  endfunction
  assign vec_data_078 = _15281_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616], data_d1[631:624] }, { _05920_, _05919_, _05918_, _05917_, _05916_, _05915_, _05914_, _05913_, _05912_, _05911_, _05910_, _05909_, _05908_, _05907_, _05906_, _05905_, _05904_, _05903_, _05902_, _05901_, _05900_, _05899_, _05898_, _05897_, _05896_, _05895_, _05894_, _05893_, _05892_, _05891_, _05890_, _05889_, _05888_, _05887_, _05886_, _05885_, _05884_, _05883_, _05882_, _05881_, _05880_, _05879_, _05878_, _05877_, _05876_, _05875_, _05874_, _05873_, _05872_, _05871_, _05870_, _05869_, _05868_, _05867_, _05866_, _05865_, _05864_, _05863_, _05862_, _05861_, _05860_, _05859_, _05858_, _05857_, _05856_, _05855_, _05854_, _05853_, _05852_, _05851_, _05850_, _05849_, _05848_, _05847_, _05846_, _05845_, _05844_, _05843_, _05842_ });
  assign _05842_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001111;
  assign _05843_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001110;
  assign _05844_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001101;
  assign _05845_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001100;
  assign _05846_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001011;
  assign _05847_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001010;
  assign _05848_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001001;
  assign _05849_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1001000;
  assign _05850_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000111;
  assign _05851_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000110;
  assign _05852_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000101;
  assign _05853_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000100;
  assign _05854_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000011;
  assign _05855_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000010;
  assign _05856_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000001;
  assign _05857_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 7'b1000000;
  assign _05858_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111111;
  assign _05859_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111110;
  assign _05860_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111101;
  assign _05861_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111100;
  assign _05862_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111011;
  assign _05863_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111010;
  assign _05864_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111001;
  assign _05865_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b111000;
  assign _05866_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110111;
  assign _05867_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110110;
  assign _05868_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110101;
  assign _05869_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110100;
  assign _05870_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110011;
  assign _05871_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110010;
  assign _05872_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110001;
  assign _05873_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b110000;
  assign _05874_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101111;
  assign _05875_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101110;
  assign _05876_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101101;
  assign _05877_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101100;
  assign _05878_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101011;
  assign _05879_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101010;
  assign _05880_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101001;
  assign _05881_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b101000;
  assign _05882_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100111;
  assign _05883_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100110;
  assign _05884_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100101;
  assign _05885_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100100;
  assign _05886_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100011;
  assign _05887_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7630|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100010;
  assign _05888_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7629|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100001;
  assign _05889_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7628|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 6'b100000;
  assign _05890_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11111;
  assign _05891_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11110;
  assign _05892_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11101;
  assign _05893_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11100;
  assign _05894_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11011;
  assign _05895_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11010;
  assign _05896_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11001;
  assign _05897_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b11000;
  assign _05898_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10111;
  assign _05899_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10110;
  assign _05900_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10101;
  assign _05901_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10100;
  assign _05902_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10011;
  assign _05903_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10010;
  assign _05904_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10001;
  assign _05905_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 5'b10000;
  assign _05906_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1111;
  assign _05907_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1110;
  assign _05908_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1101;
  assign _05909_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1100;
  assign _05910_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1011;
  assign _05911_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1010;
  assign _05912_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1001;
  assign _05913_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 4'b1000;
  assign _05914_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 3'b111;
  assign _05915_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 3'b110;
  assign _05916_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 3'b101;
  assign _05917_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 3'b100;
  assign _05918_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 2'b11;
  assign _05919_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 2'b10;
  assign _05920_ = vec_sum_078_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7596" *) 1'b1;
  function [7:0] _15361_;
    input [7:0] a;
    input [623:0] b;
    input [77:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *)
    (* parallel_case *)
    casez (s)
      78'b?????????????????????????????????????????????????????????????????????????????1:
        _15361_ = b[7:0];
      78'b????????????????????????????????????????????????????????????????????????????1?:
        _15361_ = b[15:8];
      78'b???????????????????????????????????????????????????????????????????????????1??:
        _15361_ = b[23:16];
      78'b??????????????????????????????????????????????????????????????????????????1???:
        _15361_ = b[31:24];
      78'b?????????????????????????????????????????????????????????????????????????1????:
        _15361_ = b[39:32];
      78'b????????????????????????????????????????????????????????????????????????1?????:
        _15361_ = b[47:40];
      78'b???????????????????????????????????????????????????????????????????????1??????:
        _15361_ = b[55:48];
      78'b??????????????????????????????????????????????????????????????????????1???????:
        _15361_ = b[63:56];
      78'b?????????????????????????????????????????????????????????????????????1????????:
        _15361_ = b[71:64];
      78'b????????????????????????????????????????????????????????????????????1?????????:
        _15361_ = b[79:72];
      78'b???????????????????????????????????????????????????????????????????1??????????:
        _15361_ = b[87:80];
      78'b??????????????????????????????????????????????????????????????????1???????????:
        _15361_ = b[95:88];
      78'b?????????????????????????????????????????????????????????????????1????????????:
        _15361_ = b[103:96];
      78'b????????????????????????????????????????????????????????????????1?????????????:
        _15361_ = b[111:104];
      78'b???????????????????????????????????????????????????????????????1??????????????:
        _15361_ = b[119:112];
      78'b??????????????????????????????????????????????????????????????1???????????????:
        _15361_ = b[127:120];
      78'b?????????????????????????????????????????????????????????????1????????????????:
        _15361_ = b[135:128];
      78'b????????????????????????????????????????????????????????????1?????????????????:
        _15361_ = b[143:136];
      78'b???????????????????????????????????????????????????????????1??????????????????:
        _15361_ = b[151:144];
      78'b??????????????????????????????????????????????????????????1???????????????????:
        _15361_ = b[159:152];
      78'b?????????????????????????????????????????????????????????1????????????????????:
        _15361_ = b[167:160];
      78'b????????????????????????????????????????????????????????1?????????????????????:
        _15361_ = b[175:168];
      78'b???????????????????????????????????????????????????????1??????????????????????:
        _15361_ = b[183:176];
      78'b??????????????????????????????????????????????????????1???????????????????????:
        _15361_ = b[191:184];
      78'b?????????????????????????????????????????????????????1????????????????????????:
        _15361_ = b[199:192];
      78'b????????????????????????????????????????????????????1?????????????????????????:
        _15361_ = b[207:200];
      78'b???????????????????????????????????????????????????1??????????????????????????:
        _15361_ = b[215:208];
      78'b??????????????????????????????????????????????????1???????????????????????????:
        _15361_ = b[223:216];
      78'b?????????????????????????????????????????????????1????????????????????????????:
        _15361_ = b[231:224];
      78'b????????????????????????????????????????????????1?????????????????????????????:
        _15361_ = b[239:232];
      78'b???????????????????????????????????????????????1??????????????????????????????:
        _15361_ = b[247:240];
      78'b??????????????????????????????????????????????1???????????????????????????????:
        _15361_ = b[255:248];
      78'b?????????????????????????????????????????????1????????????????????????????????:
        _15361_ = b[263:256];
      78'b????????????????????????????????????????????1?????????????????????????????????:
        _15361_ = b[271:264];
      78'b???????????????????????????????????????????1??????????????????????????????????:
        _15361_ = b[279:272];
      78'b??????????????????????????????????????????1???????????????????????????????????:
        _15361_ = b[287:280];
      78'b?????????????????????????????????????????1????????????????????????????????????:
        _15361_ = b[295:288];
      78'b????????????????????????????????????????1?????????????????????????????????????:
        _15361_ = b[303:296];
      78'b???????????????????????????????????????1??????????????????????????????????????:
        _15361_ = b[311:304];
      78'b??????????????????????????????????????1???????????????????????????????????????:
        _15361_ = b[319:312];
      78'b?????????????????????????????????????1????????????????????????????????????????:
        _15361_ = b[327:320];
      78'b????????????????????????????????????1?????????????????????????????????????????:
        _15361_ = b[335:328];
      78'b???????????????????????????????????1??????????????????????????????????????????:
        _15361_ = b[343:336];
      78'b??????????????????????????????????1???????????????????????????????????????????:
        _15361_ = b[351:344];
      78'b?????????????????????????????????1????????????????????????????????????????????:
        _15361_ = b[359:352];
      78'b????????????????????????????????1?????????????????????????????????????????????:
        _15361_ = b[367:360];
      78'b???????????????????????????????1??????????????????????????????????????????????:
        _15361_ = b[375:368];
      78'b??????????????????????????????1???????????????????????????????????????????????:
        _15361_ = b[383:376];
      78'b?????????????????????????????1????????????????????????????????????????????????:
        _15361_ = b[391:384];
      78'b????????????????????????????1?????????????????????????????????????????????????:
        _15361_ = b[399:392];
      78'b???????????????????????????1??????????????????????????????????????????????????:
        _15361_ = b[407:400];
      78'b??????????????????????????1???????????????????????????????????????????????????:
        _15361_ = b[415:408];
      78'b?????????????????????????1????????????????????????????????????????????????????:
        _15361_ = b[423:416];
      78'b????????????????????????1?????????????????????????????????????????????????????:
        _15361_ = b[431:424];
      78'b???????????????????????1??????????????????????????????????????????????????????:
        _15361_ = b[439:432];
      78'b??????????????????????1???????????????????????????????????????????????????????:
        _15361_ = b[447:440];
      78'b?????????????????????1????????????????????????????????????????????????????????:
        _15361_ = b[455:448];
      78'b????????????????????1?????????????????????????????????????????????????????????:
        _15361_ = b[463:456];
      78'b???????????????????1??????????????????????????????????????????????????????????:
        _15361_ = b[471:464];
      78'b??????????????????1???????????????????????????????????????????????????????????:
        _15361_ = b[479:472];
      78'b?????????????????1????????????????????????????????????????????????????????????:
        _15361_ = b[487:480];
      78'b????????????????1?????????????????????????????????????????????????????????????:
        _15361_ = b[495:488];
      78'b???????????????1??????????????????????????????????????????????????????????????:
        _15361_ = b[503:496];
      78'b??????????????1???????????????????????????????????????????????????????????????:
        _15361_ = b[511:504];
      78'b?????????????1????????????????????????????????????????????????????????????????:
        _15361_ = b[519:512];
      78'b????????????1?????????????????????????????????????????????????????????????????:
        _15361_ = b[527:520];
      78'b???????????1??????????????????????????????????????????????????????????????????:
        _15361_ = b[535:528];
      78'b??????????1???????????????????????????????????????????????????????????????????:
        _15361_ = b[543:536];
      78'b?????????1????????????????????????????????????????????????????????????????????:
        _15361_ = b[551:544];
      78'b????????1?????????????????????????????????????????????????????????????????????:
        _15361_ = b[559:552];
      78'b???????1??????????????????????????????????????????????????????????????????????:
        _15361_ = b[567:560];
      78'b??????1???????????????????????????????????????????????????????????????????????:
        _15361_ = b[575:568];
      78'b?????1????????????????????????????????????????????????????????????????????????:
        _15361_ = b[583:576];
      78'b????1?????????????????????????????????????????????????????????????????????????:
        _15361_ = b[591:584];
      78'b???1??????????????????????????????????????????????????????????????????????????:
        _15361_ = b[599:592];
      78'b??1???????????????????????????????????????????????????????????????????????????:
        _15361_ = b[607:600];
      78'b?1????????????????????????????????????????????????????????????????????????????:
        _15361_ = b[615:608];
      78'b1?????????????????????????????????????????????????????????????????????????????:
        _15361_ = b[623:616];
      default:
        _15361_ = a;
    endcase
  endfunction
  assign vec_data_077 = _15361_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608], data_d1[623:616] }, { _05998_, _05997_, _05996_, _05995_, _05994_, _05993_, _05992_, _05991_, _05990_, _05989_, _05988_, _05987_, _05986_, _05985_, _05984_, _05983_, _05982_, _05981_, _05980_, _05979_, _05978_, _05977_, _05976_, _05975_, _05974_, _05973_, _05972_, _05971_, _05970_, _05969_, _05968_, _05967_, _05966_, _05965_, _05964_, _05963_, _05962_, _05961_, _05960_, _05959_, _05958_, _05957_, _05956_, _05955_, _05954_, _05953_, _05952_, _05951_, _05950_, _05949_, _05948_, _05947_, _05946_, _05945_, _05944_, _05943_, _05942_, _05941_, _05940_, _05939_, _05938_, _05937_, _05936_, _05935_, _05934_, _05933_, _05932_, _05931_, _05930_, _05929_, _05928_, _05927_, _05926_, _05925_, _05924_, _05923_, _05922_, _05921_ });
  assign _05921_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001110;
  assign _05922_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001101;
  assign _05923_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001100;
  assign _05924_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001011;
  assign _05925_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001010;
  assign _05926_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001001;
  assign _05927_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1001000;
  assign _05928_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000111;
  assign _05929_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000110;
  assign _05930_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000101;
  assign _05931_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000100;
  assign _05932_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000011;
  assign _05933_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000010;
  assign _05934_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000001;
  assign _05935_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 7'b1000000;
  assign _05936_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111111;
  assign _05937_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111110;
  assign _05938_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111101;
  assign _05939_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111100;
  assign _05940_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111011;
  assign _05941_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111010;
  assign _05942_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111001;
  assign _05943_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b111000;
  assign _05944_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110111;
  assign _05945_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110110;
  assign _05946_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110101;
  assign _05947_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110100;
  assign _05948_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110011;
  assign _05949_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110010;
  assign _05950_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110001;
  assign _05951_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b110000;
  assign _05952_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101111;
  assign _05953_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101110;
  assign _05954_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101101;
  assign _05955_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101100;
  assign _05956_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101011;
  assign _05957_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101010;
  assign _05958_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101001;
  assign _05959_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b101000;
  assign _05960_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100111;
  assign _05961_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100110;
  assign _05962_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100101;
  assign _05963_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100100;
  assign _05964_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100011;
  assign _05965_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100010;
  assign _05966_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100001;
  assign _05967_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 6'b100000;
  assign _05968_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11111;
  assign _05969_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11110;
  assign _05970_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11101;
  assign _05971_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11100;
  assign _05972_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11011;
  assign _05973_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11010;
  assign _05974_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11001;
  assign _05975_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b11000;
  assign _05976_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10111;
  assign _05977_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10110;
  assign _05978_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10101;
  assign _05979_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10100;
  assign _05980_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10011;
  assign _05981_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10010;
  assign _05982_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10001;
  assign _05983_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 5'b10000;
  assign _05984_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1111;
  assign _05985_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1110;
  assign _05986_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1101;
  assign _05987_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1100;
  assign _05988_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1011;
  assign _05989_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1010;
  assign _05990_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1001;
  assign _05991_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 4'b1000;
  assign _05992_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 3'b111;
  assign _05993_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 3'b110;
  assign _05994_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 3'b101;
  assign _05995_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 3'b100;
  assign _05996_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 2'b11;
  assign _05997_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 2'b10;
  assign _05998_ = vec_sum_077_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7510" *) 1'b1;
  function [7:0] _15440_;
    input [7:0] a;
    input [615:0] b;
    input [76:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *)
    (* parallel_case *)
    casez (s)
      77'b????????????????????????????????????????????????????????????????????????????1:
        _15440_ = b[7:0];
      77'b???????????????????????????????????????????????????????????????????????????1?:
        _15440_ = b[15:8];
      77'b??????????????????????????????????????????????????????????????????????????1??:
        _15440_ = b[23:16];
      77'b?????????????????????????????????????????????????????????????????????????1???:
        _15440_ = b[31:24];
      77'b????????????????????????????????????????????????????????????????????????1????:
        _15440_ = b[39:32];
      77'b???????????????????????????????????????????????????????????????????????1?????:
        _15440_ = b[47:40];
      77'b??????????????????????????????????????????????????????????????????????1??????:
        _15440_ = b[55:48];
      77'b?????????????????????????????????????????????????????????????????????1???????:
        _15440_ = b[63:56];
      77'b????????????????????????????????????????????????????????????????????1????????:
        _15440_ = b[71:64];
      77'b???????????????????????????????????????????????????????????????????1?????????:
        _15440_ = b[79:72];
      77'b??????????????????????????????????????????????????????????????????1??????????:
        _15440_ = b[87:80];
      77'b?????????????????????????????????????????????????????????????????1???????????:
        _15440_ = b[95:88];
      77'b????????????????????????????????????????????????????????????????1????????????:
        _15440_ = b[103:96];
      77'b???????????????????????????????????????????????????????????????1?????????????:
        _15440_ = b[111:104];
      77'b??????????????????????????????????????????????????????????????1??????????????:
        _15440_ = b[119:112];
      77'b?????????????????????????????????????????????????????????????1???????????????:
        _15440_ = b[127:120];
      77'b????????????????????????????????????????????????????????????1????????????????:
        _15440_ = b[135:128];
      77'b???????????????????????????????????????????????????????????1?????????????????:
        _15440_ = b[143:136];
      77'b??????????????????????????????????????????????????????????1??????????????????:
        _15440_ = b[151:144];
      77'b?????????????????????????????????????????????????????????1???????????????????:
        _15440_ = b[159:152];
      77'b????????????????????????????????????????????????????????1????????????????????:
        _15440_ = b[167:160];
      77'b???????????????????????????????????????????????????????1?????????????????????:
        _15440_ = b[175:168];
      77'b??????????????????????????????????????????????????????1??????????????????????:
        _15440_ = b[183:176];
      77'b?????????????????????????????????????????????????????1???????????????????????:
        _15440_ = b[191:184];
      77'b????????????????????????????????????????????????????1????????????????????????:
        _15440_ = b[199:192];
      77'b???????????????????????????????????????????????????1?????????????????????????:
        _15440_ = b[207:200];
      77'b??????????????????????????????????????????????????1??????????????????????????:
        _15440_ = b[215:208];
      77'b?????????????????????????????????????????????????1???????????????????????????:
        _15440_ = b[223:216];
      77'b????????????????????????????????????????????????1????????????????????????????:
        _15440_ = b[231:224];
      77'b???????????????????????????????????????????????1?????????????????????????????:
        _15440_ = b[239:232];
      77'b??????????????????????????????????????????????1??????????????????????????????:
        _15440_ = b[247:240];
      77'b?????????????????????????????????????????????1???????????????????????????????:
        _15440_ = b[255:248];
      77'b????????????????????????????????????????????1????????????????????????????????:
        _15440_ = b[263:256];
      77'b???????????????????????????????????????????1?????????????????????????????????:
        _15440_ = b[271:264];
      77'b??????????????????????????????????????????1??????????????????????????????????:
        _15440_ = b[279:272];
      77'b?????????????????????????????????????????1???????????????????????????????????:
        _15440_ = b[287:280];
      77'b????????????????????????????????????????1????????????????????????????????????:
        _15440_ = b[295:288];
      77'b???????????????????????????????????????1?????????????????????????????????????:
        _15440_ = b[303:296];
      77'b??????????????????????????????????????1??????????????????????????????????????:
        _15440_ = b[311:304];
      77'b?????????????????????????????????????1???????????????????????????????????????:
        _15440_ = b[319:312];
      77'b????????????????????????????????????1????????????????????????????????????????:
        _15440_ = b[327:320];
      77'b???????????????????????????????????1?????????????????????????????????????????:
        _15440_ = b[335:328];
      77'b??????????????????????????????????1??????????????????????????????????????????:
        _15440_ = b[343:336];
      77'b?????????????????????????????????1???????????????????????????????????????????:
        _15440_ = b[351:344];
      77'b????????????????????????????????1????????????????????????????????????????????:
        _15440_ = b[359:352];
      77'b???????????????????????????????1?????????????????????????????????????????????:
        _15440_ = b[367:360];
      77'b??????????????????????????????1??????????????????????????????????????????????:
        _15440_ = b[375:368];
      77'b?????????????????????????????1???????????????????????????????????????????????:
        _15440_ = b[383:376];
      77'b????????????????????????????1????????????????????????????????????????????????:
        _15440_ = b[391:384];
      77'b???????????????????????????1?????????????????????????????????????????????????:
        _15440_ = b[399:392];
      77'b??????????????????????????1??????????????????????????????????????????????????:
        _15440_ = b[407:400];
      77'b?????????????????????????1???????????????????????????????????????????????????:
        _15440_ = b[415:408];
      77'b????????????????????????1????????????????????????????????????????????????????:
        _15440_ = b[423:416];
      77'b???????????????????????1?????????????????????????????????????????????????????:
        _15440_ = b[431:424];
      77'b??????????????????????1??????????????????????????????????????????????????????:
        _15440_ = b[439:432];
      77'b?????????????????????1???????????????????????????????????????????????????????:
        _15440_ = b[447:440];
      77'b????????????????????1????????????????????????????????????????????????????????:
        _15440_ = b[455:448];
      77'b???????????????????1?????????????????????????????????????????????????????????:
        _15440_ = b[463:456];
      77'b??????????????????1??????????????????????????????????????????????????????????:
        _15440_ = b[471:464];
      77'b?????????????????1???????????????????????????????????????????????????????????:
        _15440_ = b[479:472];
      77'b????????????????1????????????????????????????????????????????????????????????:
        _15440_ = b[487:480];
      77'b???????????????1?????????????????????????????????????????????????????????????:
        _15440_ = b[495:488];
      77'b??????????????1??????????????????????????????????????????????????????????????:
        _15440_ = b[503:496];
      77'b?????????????1???????????????????????????????????????????????????????????????:
        _15440_ = b[511:504];
      77'b????????????1????????????????????????????????????????????????????????????????:
        _15440_ = b[519:512];
      77'b???????????1?????????????????????????????????????????????????????????????????:
        _15440_ = b[527:520];
      77'b??????????1??????????????????????????????????????????????????????????????????:
        _15440_ = b[535:528];
      77'b?????????1???????????????????????????????????????????????????????????????????:
        _15440_ = b[543:536];
      77'b????????1????????????????????????????????????????????????????????????????????:
        _15440_ = b[551:544];
      77'b???????1?????????????????????????????????????????????????????????????????????:
        _15440_ = b[559:552];
      77'b??????1??????????????????????????????????????????????????????????????????????:
        _15440_ = b[567:560];
      77'b?????1???????????????????????????????????????????????????????????????????????:
        _15440_ = b[575:568];
      77'b????1????????????????????????????????????????????????????????????????????????:
        _15440_ = b[583:576];
      77'b???1?????????????????????????????????????????????????????????????????????????:
        _15440_ = b[591:584];
      77'b??1??????????????????????????????????????????????????????????????????????????:
        _15440_ = b[599:592];
      77'b?1???????????????????????????????????????????????????????????????????????????:
        _15440_ = b[607:600];
      77'b1????????????????????????????????????????????????????????????????????????????:
        _15440_ = b[615:608];
      default:
        _15440_ = a;
    endcase
  endfunction
  assign vec_data_076 = _15440_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600], data_d1[615:608] }, { _06075_, _06074_, _06073_, _06072_, _06071_, _06070_, _06069_, _06068_, _06067_, _06066_, _06065_, _06064_, _06063_, _06062_, _06061_, _06060_, _06059_, _06058_, _06057_, _06056_, _06055_, _06054_, _06053_, _06052_, _06051_, _06050_, _06049_, _06048_, _06047_, _06046_, _06045_, _06044_, _06043_, _06042_, _06041_, _06040_, _06039_, _06038_, _06037_, _06036_, _06035_, _06034_, _06033_, _06032_, _06031_, _06030_, _06029_, _06028_, _06027_, _06026_, _06025_, _06024_, _06023_, _06022_, _06021_, _06020_, _06019_, _06018_, _06017_, _06016_, _06015_, _06014_, _06013_, _06012_, _06011_, _06010_, _06009_, _06008_, _06007_, _06006_, _06005_, _06004_, _06003_, _06002_, _06001_, _06000_, _05999_ });
  assign _05999_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001101;
  assign _06000_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001100;
  assign _06001_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001011;
  assign _06002_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001010;
  assign _06003_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001001;
  assign _06004_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1001000;
  assign _06005_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000111;
  assign _06006_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000110;
  assign _06007_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000101;
  assign _06008_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000100;
  assign _06009_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000011;
  assign _06010_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000010;
  assign _06011_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000001;
  assign _06012_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 7'b1000000;
  assign _06013_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111111;
  assign _06014_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111110;
  assign _06015_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111101;
  assign _06016_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111100;
  assign _06017_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111011;
  assign _06018_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111010;
  assign _06019_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111001;
  assign _06020_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b111000;
  assign _06021_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110111;
  assign _06022_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110110;
  assign _06023_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110101;
  assign _06024_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110100;
  assign _06025_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110011;
  assign _06026_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110010;
  assign _06027_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110001;
  assign _06028_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b110000;
  assign _06029_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101111;
  assign _06030_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101110;
  assign _06031_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101101;
  assign _06032_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101100;
  assign _06033_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101011;
  assign _06034_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101010;
  assign _06035_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101001;
  assign _06036_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b101000;
  assign _06037_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100111;
  assign _06038_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100110;
  assign _06039_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100101;
  assign _06040_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100100;
  assign _06041_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100011;
  assign _06042_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100010;
  assign _06043_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100001;
  assign _06044_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 6'b100000;
  assign _06045_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11111;
  assign _06046_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11110;
  assign _06047_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11101;
  assign _06048_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11100;
  assign _06049_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11011;
  assign _06050_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11010;
  assign _06051_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11001;
  assign _06052_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b11000;
  assign _06053_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10111;
  assign _06054_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10110;
  assign _06055_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10101;
  assign _06056_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10100;
  assign _06057_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10011;
  assign _06058_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10010;
  assign _06059_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10001;
  assign _06060_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 5'b10000;
  assign _06061_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1111;
  assign _06062_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1110;
  assign _06063_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1101;
  assign _06064_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1100;
  assign _06065_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1011;
  assign _06066_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1010;
  assign _06067_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1001;
  assign _06068_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 4'b1000;
  assign _06069_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 3'b111;
  assign _06070_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 3'b110;
  assign _06071_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 3'b101;
  assign _06072_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 3'b100;
  assign _06073_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 2'b11;
  assign _06074_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 2'b10;
  assign _06075_ = vec_sum_076_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7425" *) 1'b1;
  function [7:0] _15518_;
    input [7:0] a;
    input [607:0] b;
    input [75:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *)
    (* parallel_case *)
    casez (s)
      76'b???????????????????????????????????????????????????????????????????????????1:
        _15518_ = b[7:0];
      76'b??????????????????????????????????????????????????????????????????????????1?:
        _15518_ = b[15:8];
      76'b?????????????????????????????????????????????????????????????????????????1??:
        _15518_ = b[23:16];
      76'b????????????????????????????????????????????????????????????????????????1???:
        _15518_ = b[31:24];
      76'b???????????????????????????????????????????????????????????????????????1????:
        _15518_ = b[39:32];
      76'b??????????????????????????????????????????????????????????????????????1?????:
        _15518_ = b[47:40];
      76'b?????????????????????????????????????????????????????????????????????1??????:
        _15518_ = b[55:48];
      76'b????????????????????????????????????????????????????????????????????1???????:
        _15518_ = b[63:56];
      76'b???????????????????????????????????????????????????????????????????1????????:
        _15518_ = b[71:64];
      76'b??????????????????????????????????????????????????????????????????1?????????:
        _15518_ = b[79:72];
      76'b?????????????????????????????????????????????????????????????????1??????????:
        _15518_ = b[87:80];
      76'b????????????????????????????????????????????????????????????????1???????????:
        _15518_ = b[95:88];
      76'b???????????????????????????????????????????????????????????????1????????????:
        _15518_ = b[103:96];
      76'b??????????????????????????????????????????????????????????????1?????????????:
        _15518_ = b[111:104];
      76'b?????????????????????????????????????????????????????????????1??????????????:
        _15518_ = b[119:112];
      76'b????????????????????????????????????????????????????????????1???????????????:
        _15518_ = b[127:120];
      76'b???????????????????????????????????????????????????????????1????????????????:
        _15518_ = b[135:128];
      76'b??????????????????????????????????????????????????????????1?????????????????:
        _15518_ = b[143:136];
      76'b?????????????????????????????????????????????????????????1??????????????????:
        _15518_ = b[151:144];
      76'b????????????????????????????????????????????????????????1???????????????????:
        _15518_ = b[159:152];
      76'b???????????????????????????????????????????????????????1????????????????????:
        _15518_ = b[167:160];
      76'b??????????????????????????????????????????????????????1?????????????????????:
        _15518_ = b[175:168];
      76'b?????????????????????????????????????????????????????1??????????????????????:
        _15518_ = b[183:176];
      76'b????????????????????????????????????????????????????1???????????????????????:
        _15518_ = b[191:184];
      76'b???????????????????????????????????????????????????1????????????????????????:
        _15518_ = b[199:192];
      76'b??????????????????????????????????????????????????1?????????????????????????:
        _15518_ = b[207:200];
      76'b?????????????????????????????????????????????????1??????????????????????????:
        _15518_ = b[215:208];
      76'b????????????????????????????????????????????????1???????????????????????????:
        _15518_ = b[223:216];
      76'b???????????????????????????????????????????????1????????????????????????????:
        _15518_ = b[231:224];
      76'b??????????????????????????????????????????????1?????????????????????????????:
        _15518_ = b[239:232];
      76'b?????????????????????????????????????????????1??????????????????????????????:
        _15518_ = b[247:240];
      76'b????????????????????????????????????????????1???????????????????????????????:
        _15518_ = b[255:248];
      76'b???????????????????????????????????????????1????????????????????????????????:
        _15518_ = b[263:256];
      76'b??????????????????????????????????????????1?????????????????????????????????:
        _15518_ = b[271:264];
      76'b?????????????????????????????????????????1??????????????????????????????????:
        _15518_ = b[279:272];
      76'b????????????????????????????????????????1???????????????????????????????????:
        _15518_ = b[287:280];
      76'b???????????????????????????????????????1????????????????????????????????????:
        _15518_ = b[295:288];
      76'b??????????????????????????????????????1?????????????????????????????????????:
        _15518_ = b[303:296];
      76'b?????????????????????????????????????1??????????????????????????????????????:
        _15518_ = b[311:304];
      76'b????????????????????????????????????1???????????????????????????????????????:
        _15518_ = b[319:312];
      76'b???????????????????????????????????1????????????????????????????????????????:
        _15518_ = b[327:320];
      76'b??????????????????????????????????1?????????????????????????????????????????:
        _15518_ = b[335:328];
      76'b?????????????????????????????????1??????????????????????????????????????????:
        _15518_ = b[343:336];
      76'b????????????????????????????????1???????????????????????????????????????????:
        _15518_ = b[351:344];
      76'b???????????????????????????????1????????????????????????????????????????????:
        _15518_ = b[359:352];
      76'b??????????????????????????????1?????????????????????????????????????????????:
        _15518_ = b[367:360];
      76'b?????????????????????????????1??????????????????????????????????????????????:
        _15518_ = b[375:368];
      76'b????????????????????????????1???????????????????????????????????????????????:
        _15518_ = b[383:376];
      76'b???????????????????????????1????????????????????????????????????????????????:
        _15518_ = b[391:384];
      76'b??????????????????????????1?????????????????????????????????????????????????:
        _15518_ = b[399:392];
      76'b?????????????????????????1??????????????????????????????????????????????????:
        _15518_ = b[407:400];
      76'b????????????????????????1???????????????????????????????????????????????????:
        _15518_ = b[415:408];
      76'b???????????????????????1????????????????????????????????????????????????????:
        _15518_ = b[423:416];
      76'b??????????????????????1?????????????????????????????????????????????????????:
        _15518_ = b[431:424];
      76'b?????????????????????1??????????????????????????????????????????????????????:
        _15518_ = b[439:432];
      76'b????????????????????1???????????????????????????????????????????????????????:
        _15518_ = b[447:440];
      76'b???????????????????1????????????????????????????????????????????????????????:
        _15518_ = b[455:448];
      76'b??????????????????1?????????????????????????????????????????????????????????:
        _15518_ = b[463:456];
      76'b?????????????????1??????????????????????????????????????????????????????????:
        _15518_ = b[471:464];
      76'b????????????????1???????????????????????????????????????????????????????????:
        _15518_ = b[479:472];
      76'b???????????????1????????????????????????????????????????????????????????????:
        _15518_ = b[487:480];
      76'b??????????????1?????????????????????????????????????????????????????????????:
        _15518_ = b[495:488];
      76'b?????????????1??????????????????????????????????????????????????????????????:
        _15518_ = b[503:496];
      76'b????????????1???????????????????????????????????????????????????????????????:
        _15518_ = b[511:504];
      76'b???????????1????????????????????????????????????????????????????????????????:
        _15518_ = b[519:512];
      76'b??????????1?????????????????????????????????????????????????????????????????:
        _15518_ = b[527:520];
      76'b?????????1??????????????????????????????????????????????????????????????????:
        _15518_ = b[535:528];
      76'b????????1???????????????????????????????????????????????????????????????????:
        _15518_ = b[543:536];
      76'b???????1????????????????????????????????????????????????????????????????????:
        _15518_ = b[551:544];
      76'b??????1?????????????????????????????????????????????????????????????????????:
        _15518_ = b[559:552];
      76'b?????1??????????????????????????????????????????????????????????????????????:
        _15518_ = b[567:560];
      76'b????1???????????????????????????????????????????????????????????????????????:
        _15518_ = b[575:568];
      76'b???1????????????????????????????????????????????????????????????????????????:
        _15518_ = b[583:576];
      76'b??1?????????????????????????????????????????????????????????????????????????:
        _15518_ = b[591:584];
      76'b?1??????????????????????????????????????????????????????????????????????????:
        _15518_ = b[599:592];
      76'b1???????????????????????????????????????????????????????????????????????????:
        _15518_ = b[607:600];
      default:
        _15518_ = a;
    endcase
  endfunction
  assign vec_data_075 = _15518_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592], data_d1[607:600] }, { _06151_, _06150_, _06149_, _06148_, _06147_, _06146_, _06145_, _06144_, _06143_, _06142_, _06141_, _06140_, _06139_, _06138_, _06137_, _06136_, _06135_, _06134_, _06133_, _06132_, _06131_, _06130_, _06129_, _06128_, _06127_, _06126_, _06125_, _06124_, _06123_, _06122_, _06121_, _06120_, _06119_, _06118_, _06117_, _06116_, _06115_, _06114_, _06113_, _06112_, _06111_, _06110_, _06109_, _06108_, _06107_, _06106_, _06105_, _06104_, _06103_, _06102_, _06101_, _06100_, _06099_, _06098_, _06097_, _06096_, _06095_, _06094_, _06093_, _06092_, _06091_, _06090_, _06089_, _06088_, _06087_, _06086_, _06085_, _06084_, _06083_, _06082_, _06081_, _06080_, _06079_, _06078_, _06077_, _06076_ });
  assign _06076_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1001100;
  assign _06077_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1001011;
  assign _06078_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1001010;
  assign _06079_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1001001;
  assign _06080_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1001000;
  assign _06081_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000111;
  assign _06082_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000110;
  assign _06083_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7410|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000101;
  assign _06084_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7409|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000100;
  assign _06085_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000011;
  assign _06086_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000010;
  assign _06087_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000001;
  assign _06088_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 7'b1000000;
  assign _06089_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111111;
  assign _06090_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111110;
  assign _06091_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111101;
  assign _06092_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111100;
  assign _06093_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111011;
  assign _06094_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111010;
  assign _06095_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111001;
  assign _06096_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b111000;
  assign _06097_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110111;
  assign _06098_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110110;
  assign _06099_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110101;
  assign _06100_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110100;
  assign _06101_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110011;
  assign _06102_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110010;
  assign _06103_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110001;
  assign _06104_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b110000;
  assign _06105_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101111;
  assign _06106_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101110;
  assign _06107_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101101;
  assign _06108_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101100;
  assign _06109_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101011;
  assign _06110_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101010;
  assign _06111_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101001;
  assign _06112_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b101000;
  assign _06113_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100111;
  assign _06114_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100110;
  assign _06115_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100101;
  assign _06116_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100100;
  assign _06117_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100011;
  assign _06118_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100010;
  assign _06119_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100001;
  assign _06120_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 6'b100000;
  assign _06121_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11111;
  assign _06122_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11110;
  assign _06123_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11101;
  assign _06124_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11100;
  assign _06125_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11011;
  assign _06126_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11010;
  assign _06127_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11001;
  assign _06128_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b11000;
  assign _06129_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10111;
  assign _06130_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10110;
  assign _06131_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10101;
  assign _06132_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10100;
  assign _06133_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10011;
  assign _06134_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10010;
  assign _06135_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10001;
  assign _06136_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 5'b10000;
  assign _06137_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1111;
  assign _06138_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1110;
  assign _06139_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1101;
  assign _06140_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1100;
  assign _06141_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1011;
  assign _06142_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1010;
  assign _06143_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1001;
  assign _06144_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 4'b1000;
  assign _06145_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 3'b111;
  assign _06146_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 3'b110;
  assign _06147_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 3'b101;
  assign _06148_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 3'b100;
  assign _06149_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 2'b11;
  assign _06150_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 2'b10;
  assign _06151_ = vec_sum_075_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7341" *) 1'b1;
  function [7:0] _15595_;
    input [7:0] a;
    input [599:0] b;
    input [74:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *)
    (* parallel_case *)
    casez (s)
      75'b??????????????????????????????????????????????????????????????????????????1:
        _15595_ = b[7:0];
      75'b?????????????????????????????????????????????????????????????????????????1?:
        _15595_ = b[15:8];
      75'b????????????????????????????????????????????????????????????????????????1??:
        _15595_ = b[23:16];
      75'b???????????????????????????????????????????????????????????????????????1???:
        _15595_ = b[31:24];
      75'b??????????????????????????????????????????????????????????????????????1????:
        _15595_ = b[39:32];
      75'b?????????????????????????????????????????????????????????????????????1?????:
        _15595_ = b[47:40];
      75'b????????????????????????????????????????????????????????????????????1??????:
        _15595_ = b[55:48];
      75'b???????????????????????????????????????????????????????????????????1???????:
        _15595_ = b[63:56];
      75'b??????????????????????????????????????????????????????????????????1????????:
        _15595_ = b[71:64];
      75'b?????????????????????????????????????????????????????????????????1?????????:
        _15595_ = b[79:72];
      75'b????????????????????????????????????????????????????????????????1??????????:
        _15595_ = b[87:80];
      75'b???????????????????????????????????????????????????????????????1???????????:
        _15595_ = b[95:88];
      75'b??????????????????????????????????????????????????????????????1????????????:
        _15595_ = b[103:96];
      75'b?????????????????????????????????????????????????????????????1?????????????:
        _15595_ = b[111:104];
      75'b????????????????????????????????????????????????????????????1??????????????:
        _15595_ = b[119:112];
      75'b???????????????????????????????????????????????????????????1???????????????:
        _15595_ = b[127:120];
      75'b??????????????????????????????????????????????????????????1????????????????:
        _15595_ = b[135:128];
      75'b?????????????????????????????????????????????????????????1?????????????????:
        _15595_ = b[143:136];
      75'b????????????????????????????????????????????????????????1??????????????????:
        _15595_ = b[151:144];
      75'b???????????????????????????????????????????????????????1???????????????????:
        _15595_ = b[159:152];
      75'b??????????????????????????????????????????????????????1????????????????????:
        _15595_ = b[167:160];
      75'b?????????????????????????????????????????????????????1?????????????????????:
        _15595_ = b[175:168];
      75'b????????????????????????????????????????????????????1??????????????????????:
        _15595_ = b[183:176];
      75'b???????????????????????????????????????????????????1???????????????????????:
        _15595_ = b[191:184];
      75'b??????????????????????????????????????????????????1????????????????????????:
        _15595_ = b[199:192];
      75'b?????????????????????????????????????????????????1?????????????????????????:
        _15595_ = b[207:200];
      75'b????????????????????????????????????????????????1??????????????????????????:
        _15595_ = b[215:208];
      75'b???????????????????????????????????????????????1???????????????????????????:
        _15595_ = b[223:216];
      75'b??????????????????????????????????????????????1????????????????????????????:
        _15595_ = b[231:224];
      75'b?????????????????????????????????????????????1?????????????????????????????:
        _15595_ = b[239:232];
      75'b????????????????????????????????????????????1??????????????????????????????:
        _15595_ = b[247:240];
      75'b???????????????????????????????????????????1???????????????????????????????:
        _15595_ = b[255:248];
      75'b??????????????????????????????????????????1????????????????????????????????:
        _15595_ = b[263:256];
      75'b?????????????????????????????????????????1?????????????????????????????????:
        _15595_ = b[271:264];
      75'b????????????????????????????????????????1??????????????????????????????????:
        _15595_ = b[279:272];
      75'b???????????????????????????????????????1???????????????????????????????????:
        _15595_ = b[287:280];
      75'b??????????????????????????????????????1????????????????????????????????????:
        _15595_ = b[295:288];
      75'b?????????????????????????????????????1?????????????????????????????????????:
        _15595_ = b[303:296];
      75'b????????????????????????????????????1??????????????????????????????????????:
        _15595_ = b[311:304];
      75'b???????????????????????????????????1???????????????????????????????????????:
        _15595_ = b[319:312];
      75'b??????????????????????????????????1????????????????????????????????????????:
        _15595_ = b[327:320];
      75'b?????????????????????????????????1?????????????????????????????????????????:
        _15595_ = b[335:328];
      75'b????????????????????????????????1??????????????????????????????????????????:
        _15595_ = b[343:336];
      75'b???????????????????????????????1???????????????????????????????????????????:
        _15595_ = b[351:344];
      75'b??????????????????????????????1????????????????????????????????????????????:
        _15595_ = b[359:352];
      75'b?????????????????????????????1?????????????????????????????????????????????:
        _15595_ = b[367:360];
      75'b????????????????????????????1??????????????????????????????????????????????:
        _15595_ = b[375:368];
      75'b???????????????????????????1???????????????????????????????????????????????:
        _15595_ = b[383:376];
      75'b??????????????????????????1????????????????????????????????????????????????:
        _15595_ = b[391:384];
      75'b?????????????????????????1?????????????????????????????????????????????????:
        _15595_ = b[399:392];
      75'b????????????????????????1??????????????????????????????????????????????????:
        _15595_ = b[407:400];
      75'b???????????????????????1???????????????????????????????????????????????????:
        _15595_ = b[415:408];
      75'b??????????????????????1????????????????????????????????????????????????????:
        _15595_ = b[423:416];
      75'b?????????????????????1?????????????????????????????????????????????????????:
        _15595_ = b[431:424];
      75'b????????????????????1??????????????????????????????????????????????????????:
        _15595_ = b[439:432];
      75'b???????????????????1???????????????????????????????????????????????????????:
        _15595_ = b[447:440];
      75'b??????????????????1????????????????????????????????????????????????????????:
        _15595_ = b[455:448];
      75'b?????????????????1?????????????????????????????????????????????????????????:
        _15595_ = b[463:456];
      75'b????????????????1??????????????????????????????????????????????????????????:
        _15595_ = b[471:464];
      75'b???????????????1???????????????????????????????????????????????????????????:
        _15595_ = b[479:472];
      75'b??????????????1????????????????????????????????????????????????????????????:
        _15595_ = b[487:480];
      75'b?????????????1?????????????????????????????????????????????????????????????:
        _15595_ = b[495:488];
      75'b????????????1??????????????????????????????????????????????????????????????:
        _15595_ = b[503:496];
      75'b???????????1???????????????????????????????????????????????????????????????:
        _15595_ = b[511:504];
      75'b??????????1????????????????????????????????????????????????????????????????:
        _15595_ = b[519:512];
      75'b?????????1?????????????????????????????????????????????????????????????????:
        _15595_ = b[527:520];
      75'b????????1??????????????????????????????????????????????????????????????????:
        _15595_ = b[535:528];
      75'b???????1???????????????????????????????????????????????????????????????????:
        _15595_ = b[543:536];
      75'b??????1????????????????????????????????????????????????????????????????????:
        _15595_ = b[551:544];
      75'b?????1?????????????????????????????????????????????????????????????????????:
        _15595_ = b[559:552];
      75'b????1??????????????????????????????????????????????????????????????????????:
        _15595_ = b[567:560];
      75'b???1???????????????????????????????????????????????????????????????????????:
        _15595_ = b[575:568];
      75'b??1????????????????????????????????????????????????????????????????????????:
        _15595_ = b[583:576];
      75'b?1?????????????????????????????????????????????????????????????????????????:
        _15595_ = b[591:584];
      75'b1??????????????????????????????????????????????????????????????????????????:
        _15595_ = b[599:592];
      default:
        _15595_ = a;
    endcase
  endfunction
  assign vec_data_074 = _15595_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584], data_d1[599:592] }, { _06226_, _06225_, _06224_, _06223_, _06222_, _06221_, _06220_, _06219_, _06218_, _06217_, _06216_, _06215_, _06214_, _06213_, _06212_, _06211_, _06210_, _06209_, _06208_, _06207_, _06206_, _06205_, _06204_, _06203_, _06202_, _06201_, _06200_, _06199_, _06198_, _06197_, _06196_, _06195_, _06194_, _06193_, _06192_, _06191_, _06190_, _06189_, _06188_, _06187_, _06186_, _06185_, _06184_, _06183_, _06182_, _06181_, _06180_, _06179_, _06178_, _06177_, _06176_, _06175_, _06174_, _06173_, _06172_, _06171_, _06170_, _06169_, _06168_, _06167_, _06166_, _06165_, _06164_, _06163_, _06162_, _06161_, _06160_, _06159_, _06158_, _06157_, _06156_, _06155_, _06154_, _06153_, _06152_ });
  assign _06152_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1001011;
  assign _06153_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1001010;
  assign _06154_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1001001;
  assign _06155_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1001000;
  assign _06156_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000111;
  assign _06157_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000110;
  assign _06158_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000101;
  assign _06159_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000100;
  assign _06160_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000011;
  assign _06161_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000010;
  assign _06162_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000001;
  assign _06163_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 7'b1000000;
  assign _06164_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111111;
  assign _06165_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111110;
  assign _06166_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111101;
  assign _06167_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111100;
  assign _06168_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111011;
  assign _06169_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111010;
  assign _06170_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111001;
  assign _06171_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b111000;
  assign _06172_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110111;
  assign _06173_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110110;
  assign _06174_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110101;
  assign _06175_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110100;
  assign _06176_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110011;
  assign _06177_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110010;
  assign _06178_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110001;
  assign _06179_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b110000;
  assign _06180_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101111;
  assign _06181_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101110;
  assign _06182_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101101;
  assign _06183_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101100;
  assign _06184_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101011;
  assign _06185_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101010;
  assign _06186_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101001;
  assign _06187_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b101000;
  assign _06188_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100111;
  assign _06189_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100110;
  assign _06190_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100101;
  assign _06191_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100100;
  assign _06192_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100011;
  assign _06193_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100010;
  assign _06194_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100001;
  assign _06195_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 6'b100000;
  assign _06196_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11111;
  assign _06197_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11110;
  assign _06198_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11101;
  assign _06199_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11100;
  assign _06200_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11011;
  assign _06201_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11010;
  assign _06202_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11001;
  assign _06203_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b11000;
  assign _06204_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10111;
  assign _06205_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10110;
  assign _06206_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10101;
  assign _06207_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10100;
  assign _06208_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10011;
  assign _06209_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10010;
  assign _06210_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10001;
  assign _06211_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 5'b10000;
  assign _06212_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1111;
  assign _06213_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1110;
  assign _06214_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1101;
  assign _06215_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1100;
  assign _06216_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1011;
  assign _06217_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1010;
  assign _06218_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1001;
  assign _06219_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 4'b1000;
  assign _06220_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 3'b111;
  assign _06221_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 3'b110;
  assign _06222_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 3'b101;
  assign _06223_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 3'b100;
  assign _06224_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 2'b11;
  assign _06225_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 2'b10;
  assign _06226_ = vec_sum_074_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7258" *) 1'b1;
  function [7:0] _15671_;
    input [7:0] a;
    input [591:0] b;
    input [73:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *)
    (* parallel_case *)
    casez (s)
      74'b?????????????????????????????????????????????????????????????????????????1:
        _15671_ = b[7:0];
      74'b????????????????????????????????????????????????????????????????????????1?:
        _15671_ = b[15:8];
      74'b???????????????????????????????????????????????????????????????????????1??:
        _15671_ = b[23:16];
      74'b??????????????????????????????????????????????????????????????????????1???:
        _15671_ = b[31:24];
      74'b?????????????????????????????????????????????????????????????????????1????:
        _15671_ = b[39:32];
      74'b????????????????????????????????????????????????????????????????????1?????:
        _15671_ = b[47:40];
      74'b???????????????????????????????????????????????????????????????????1??????:
        _15671_ = b[55:48];
      74'b??????????????????????????????????????????????????????????????????1???????:
        _15671_ = b[63:56];
      74'b?????????????????????????????????????????????????????????????????1????????:
        _15671_ = b[71:64];
      74'b????????????????????????????????????????????????????????????????1?????????:
        _15671_ = b[79:72];
      74'b???????????????????????????????????????????????????????????????1??????????:
        _15671_ = b[87:80];
      74'b??????????????????????????????????????????????????????????????1???????????:
        _15671_ = b[95:88];
      74'b?????????????????????????????????????????????????????????????1????????????:
        _15671_ = b[103:96];
      74'b????????????????????????????????????????????????????????????1?????????????:
        _15671_ = b[111:104];
      74'b???????????????????????????????????????????????????????????1??????????????:
        _15671_ = b[119:112];
      74'b??????????????????????????????????????????????????????????1???????????????:
        _15671_ = b[127:120];
      74'b?????????????????????????????????????????????????????????1????????????????:
        _15671_ = b[135:128];
      74'b????????????????????????????????????????????????????????1?????????????????:
        _15671_ = b[143:136];
      74'b???????????????????????????????????????????????????????1??????????????????:
        _15671_ = b[151:144];
      74'b??????????????????????????????????????????????????????1???????????????????:
        _15671_ = b[159:152];
      74'b?????????????????????????????????????????????????????1????????????????????:
        _15671_ = b[167:160];
      74'b????????????????????????????????????????????????????1?????????????????????:
        _15671_ = b[175:168];
      74'b???????????????????????????????????????????????????1??????????????????????:
        _15671_ = b[183:176];
      74'b??????????????????????????????????????????????????1???????????????????????:
        _15671_ = b[191:184];
      74'b?????????????????????????????????????????????????1????????????????????????:
        _15671_ = b[199:192];
      74'b????????????????????????????????????????????????1?????????????????????????:
        _15671_ = b[207:200];
      74'b???????????????????????????????????????????????1??????????????????????????:
        _15671_ = b[215:208];
      74'b??????????????????????????????????????????????1???????????????????????????:
        _15671_ = b[223:216];
      74'b?????????????????????????????????????????????1????????????????????????????:
        _15671_ = b[231:224];
      74'b????????????????????????????????????????????1?????????????????????????????:
        _15671_ = b[239:232];
      74'b???????????????????????????????????????????1??????????????????????????????:
        _15671_ = b[247:240];
      74'b??????????????????????????????????????????1???????????????????????????????:
        _15671_ = b[255:248];
      74'b?????????????????????????????????????????1????????????????????????????????:
        _15671_ = b[263:256];
      74'b????????????????????????????????????????1?????????????????????????????????:
        _15671_ = b[271:264];
      74'b???????????????????????????????????????1??????????????????????????????????:
        _15671_ = b[279:272];
      74'b??????????????????????????????????????1???????????????????????????????????:
        _15671_ = b[287:280];
      74'b?????????????????????????????????????1????????????????????????????????????:
        _15671_ = b[295:288];
      74'b????????????????????????????????????1?????????????????????????????????????:
        _15671_ = b[303:296];
      74'b???????????????????????????????????1??????????????????????????????????????:
        _15671_ = b[311:304];
      74'b??????????????????????????????????1???????????????????????????????????????:
        _15671_ = b[319:312];
      74'b?????????????????????????????????1????????????????????????????????????????:
        _15671_ = b[327:320];
      74'b????????????????????????????????1?????????????????????????????????????????:
        _15671_ = b[335:328];
      74'b???????????????????????????????1??????????????????????????????????????????:
        _15671_ = b[343:336];
      74'b??????????????????????????????1???????????????????????????????????????????:
        _15671_ = b[351:344];
      74'b?????????????????????????????1????????????????????????????????????????????:
        _15671_ = b[359:352];
      74'b????????????????????????????1?????????????????????????????????????????????:
        _15671_ = b[367:360];
      74'b???????????????????????????1??????????????????????????????????????????????:
        _15671_ = b[375:368];
      74'b??????????????????????????1???????????????????????????????????????????????:
        _15671_ = b[383:376];
      74'b?????????????????????????1????????????????????????????????????????????????:
        _15671_ = b[391:384];
      74'b????????????????????????1?????????????????????????????????????????????????:
        _15671_ = b[399:392];
      74'b???????????????????????1??????????????????????????????????????????????????:
        _15671_ = b[407:400];
      74'b??????????????????????1???????????????????????????????????????????????????:
        _15671_ = b[415:408];
      74'b?????????????????????1????????????????????????????????????????????????????:
        _15671_ = b[423:416];
      74'b????????????????????1?????????????????????????????????????????????????????:
        _15671_ = b[431:424];
      74'b???????????????????1??????????????????????????????????????????????????????:
        _15671_ = b[439:432];
      74'b??????????????????1???????????????????????????????????????????????????????:
        _15671_ = b[447:440];
      74'b?????????????????1????????????????????????????????????????????????????????:
        _15671_ = b[455:448];
      74'b????????????????1?????????????????????????????????????????????????????????:
        _15671_ = b[463:456];
      74'b???????????????1??????????????????????????????????????????????????????????:
        _15671_ = b[471:464];
      74'b??????????????1???????????????????????????????????????????????????????????:
        _15671_ = b[479:472];
      74'b?????????????1????????????????????????????????????????????????????????????:
        _15671_ = b[487:480];
      74'b????????????1?????????????????????????????????????????????????????????????:
        _15671_ = b[495:488];
      74'b???????????1??????????????????????????????????????????????????????????????:
        _15671_ = b[503:496];
      74'b??????????1???????????????????????????????????????????????????????????????:
        _15671_ = b[511:504];
      74'b?????????1????????????????????????????????????????????????????????????????:
        _15671_ = b[519:512];
      74'b????????1?????????????????????????????????????????????????????????????????:
        _15671_ = b[527:520];
      74'b???????1??????????????????????????????????????????????????????????????????:
        _15671_ = b[535:528];
      74'b??????1???????????????????????????????????????????????????????????????????:
        _15671_ = b[543:536];
      74'b?????1????????????????????????????????????????????????????????????????????:
        _15671_ = b[551:544];
      74'b????1?????????????????????????????????????????????????????????????????????:
        _15671_ = b[559:552];
      74'b???1??????????????????????????????????????????????????????????????????????:
        _15671_ = b[567:560];
      74'b??1???????????????????????????????????????????????????????????????????????:
        _15671_ = b[575:568];
      74'b?1????????????????????????????????????????????????????????????????????????:
        _15671_ = b[583:576];
      74'b1?????????????????????????????????????????????????????????????????????????:
        _15671_ = b[591:584];
      default:
        _15671_ = a;
    endcase
  endfunction
  assign vec_data_073 = _15671_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576], data_d1[591:584] }, { _06300_, _06299_, _06298_, _06297_, _06296_, _06295_, _06294_, _06293_, _06292_, _06291_, _06290_, _06289_, _06288_, _06287_, _06286_, _06285_, _06284_, _06283_, _06282_, _06281_, _06280_, _06279_, _06278_, _06277_, _06276_, _06275_, _06274_, _06273_, _06272_, _06271_, _06270_, _06269_, _06268_, _06267_, _06266_, _06265_, _06264_, _06263_, _06262_, _06261_, _06260_, _06259_, _06258_, _06257_, _06256_, _06255_, _06254_, _06253_, _06252_, _06251_, _06250_, _06249_, _06248_, _06247_, _06246_, _06245_, _06244_, _06243_, _06242_, _06241_, _06240_, _06239_, _06238_, _06237_, _06236_, _06235_, _06234_, _06233_, _06232_, _06231_, _06230_, _06229_, _06228_, _06227_ });
  assign _06227_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1001010;
  assign _06228_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1001001;
  assign _06229_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1001000;
  assign _06230_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000111;
  assign _06231_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000110;
  assign _06232_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000101;
  assign _06233_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000100;
  assign _06234_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000011;
  assign _06235_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000010;
  assign _06236_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000001;
  assign _06237_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 7'b1000000;
  assign _06238_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111111;
  assign _06239_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111110;
  assign _06240_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111101;
  assign _06241_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111100;
  assign _06242_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111011;
  assign _06243_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111010;
  assign _06244_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7233|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111001;
  assign _06245_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b111000;
  assign _06246_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110111;
  assign _06247_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110110;
  assign _06248_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110101;
  assign _06249_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110100;
  assign _06250_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110011;
  assign _06251_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110010;
  assign _06252_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110001;
  assign _06253_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b110000;
  assign _06254_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101111;
  assign _06255_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101110;
  assign _06256_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101101;
  assign _06257_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101100;
  assign _06258_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101011;
  assign _06259_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101010;
  assign _06260_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101001;
  assign _06261_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b101000;
  assign _06262_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100111;
  assign _06263_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100110;
  assign _06264_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100101;
  assign _06265_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100100;
  assign _06266_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100011;
  assign _06267_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100010;
  assign _06268_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100001;
  assign _06269_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 6'b100000;
  assign _06270_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11111;
  assign _06271_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11110;
  assign _06272_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11101;
  assign _06273_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11100;
  assign _06274_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11011;
  assign _06275_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11010;
  assign _06276_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11001;
  assign _06277_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b11000;
  assign _06278_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10111;
  assign _06279_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10110;
  assign _06280_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10101;
  assign _06281_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10100;
  assign _06282_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10011;
  assign _06283_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10010;
  assign _06284_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10001;
  assign _06285_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 5'b10000;
  assign _06286_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1111;
  assign _06287_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1110;
  assign _06288_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1101;
  assign _06289_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1100;
  assign _06290_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1011;
  assign _06291_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1010;
  assign _06292_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1001;
  assign _06293_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 4'b1000;
  assign _06294_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 3'b111;
  assign _06295_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 3'b110;
  assign _06296_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 3'b101;
  assign _06297_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 3'b100;
  assign _06298_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 2'b11;
  assign _06299_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 2'b10;
  assign _06300_ = vec_sum_073_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7176" *) 1'b1;
  function [7:0] _15746_;
    input [7:0] a;
    input [583:0] b;
    input [72:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *)
    (* parallel_case *)
    casez (s)
      73'b????????????????????????????????????????????????????????????????????????1:
        _15746_ = b[7:0];
      73'b???????????????????????????????????????????????????????????????????????1?:
        _15746_ = b[15:8];
      73'b??????????????????????????????????????????????????????????????????????1??:
        _15746_ = b[23:16];
      73'b?????????????????????????????????????????????????????????????????????1???:
        _15746_ = b[31:24];
      73'b????????????????????????????????????????????????????????????????????1????:
        _15746_ = b[39:32];
      73'b???????????????????????????????????????????????????????????????????1?????:
        _15746_ = b[47:40];
      73'b??????????????????????????????????????????????????????????????????1??????:
        _15746_ = b[55:48];
      73'b?????????????????????????????????????????????????????????????????1???????:
        _15746_ = b[63:56];
      73'b????????????????????????????????????????????????????????????????1????????:
        _15746_ = b[71:64];
      73'b???????????????????????????????????????????????????????????????1?????????:
        _15746_ = b[79:72];
      73'b??????????????????????????????????????????????????????????????1??????????:
        _15746_ = b[87:80];
      73'b?????????????????????????????????????????????????????????????1???????????:
        _15746_ = b[95:88];
      73'b????????????????????????????????????????????????????????????1????????????:
        _15746_ = b[103:96];
      73'b???????????????????????????????????????????????????????????1?????????????:
        _15746_ = b[111:104];
      73'b??????????????????????????????????????????????????????????1??????????????:
        _15746_ = b[119:112];
      73'b?????????????????????????????????????????????????????????1???????????????:
        _15746_ = b[127:120];
      73'b????????????????????????????????????????????????????????1????????????????:
        _15746_ = b[135:128];
      73'b???????????????????????????????????????????????????????1?????????????????:
        _15746_ = b[143:136];
      73'b??????????????????????????????????????????????????????1??????????????????:
        _15746_ = b[151:144];
      73'b?????????????????????????????????????????????????????1???????????????????:
        _15746_ = b[159:152];
      73'b????????????????????????????????????????????????????1????????????????????:
        _15746_ = b[167:160];
      73'b???????????????????????????????????????????????????1?????????????????????:
        _15746_ = b[175:168];
      73'b??????????????????????????????????????????????????1??????????????????????:
        _15746_ = b[183:176];
      73'b?????????????????????????????????????????????????1???????????????????????:
        _15746_ = b[191:184];
      73'b????????????????????????????????????????????????1????????????????????????:
        _15746_ = b[199:192];
      73'b???????????????????????????????????????????????1?????????????????????????:
        _15746_ = b[207:200];
      73'b??????????????????????????????????????????????1??????????????????????????:
        _15746_ = b[215:208];
      73'b?????????????????????????????????????????????1???????????????????????????:
        _15746_ = b[223:216];
      73'b????????????????????????????????????????????1????????????????????????????:
        _15746_ = b[231:224];
      73'b???????????????????????????????????????????1?????????????????????????????:
        _15746_ = b[239:232];
      73'b??????????????????????????????????????????1??????????????????????????????:
        _15746_ = b[247:240];
      73'b?????????????????????????????????????????1???????????????????????????????:
        _15746_ = b[255:248];
      73'b????????????????????????????????????????1????????????????????????????????:
        _15746_ = b[263:256];
      73'b???????????????????????????????????????1?????????????????????????????????:
        _15746_ = b[271:264];
      73'b??????????????????????????????????????1??????????????????????????????????:
        _15746_ = b[279:272];
      73'b?????????????????????????????????????1???????????????????????????????????:
        _15746_ = b[287:280];
      73'b????????????????????????????????????1????????????????????????????????????:
        _15746_ = b[295:288];
      73'b???????????????????????????????????1?????????????????????????????????????:
        _15746_ = b[303:296];
      73'b??????????????????????????????????1??????????????????????????????????????:
        _15746_ = b[311:304];
      73'b?????????????????????????????????1???????????????????????????????????????:
        _15746_ = b[319:312];
      73'b????????????????????????????????1????????????????????????????????????????:
        _15746_ = b[327:320];
      73'b???????????????????????????????1?????????????????????????????????????????:
        _15746_ = b[335:328];
      73'b??????????????????????????????1??????????????????????????????????????????:
        _15746_ = b[343:336];
      73'b?????????????????????????????1???????????????????????????????????????????:
        _15746_ = b[351:344];
      73'b????????????????????????????1????????????????????????????????????????????:
        _15746_ = b[359:352];
      73'b???????????????????????????1?????????????????????????????????????????????:
        _15746_ = b[367:360];
      73'b??????????????????????????1??????????????????????????????????????????????:
        _15746_ = b[375:368];
      73'b?????????????????????????1???????????????????????????????????????????????:
        _15746_ = b[383:376];
      73'b????????????????????????1????????????????????????????????????????????????:
        _15746_ = b[391:384];
      73'b???????????????????????1?????????????????????????????????????????????????:
        _15746_ = b[399:392];
      73'b??????????????????????1??????????????????????????????????????????????????:
        _15746_ = b[407:400];
      73'b?????????????????????1???????????????????????????????????????????????????:
        _15746_ = b[415:408];
      73'b????????????????????1????????????????????????????????????????????????????:
        _15746_ = b[423:416];
      73'b???????????????????1?????????????????????????????????????????????????????:
        _15746_ = b[431:424];
      73'b??????????????????1??????????????????????????????????????????????????????:
        _15746_ = b[439:432];
      73'b?????????????????1???????????????????????????????????????????????????????:
        _15746_ = b[447:440];
      73'b????????????????1????????????????????????????????????????????????????????:
        _15746_ = b[455:448];
      73'b???????????????1?????????????????????????????????????????????????????????:
        _15746_ = b[463:456];
      73'b??????????????1??????????????????????????????????????????????????????????:
        _15746_ = b[471:464];
      73'b?????????????1???????????????????????????????????????????????????????????:
        _15746_ = b[479:472];
      73'b????????????1????????????????????????????????????????????????????????????:
        _15746_ = b[487:480];
      73'b???????????1?????????????????????????????????????????????????????????????:
        _15746_ = b[495:488];
      73'b??????????1??????????????????????????????????????????????????????????????:
        _15746_ = b[503:496];
      73'b?????????1???????????????????????????????????????????????????????????????:
        _15746_ = b[511:504];
      73'b????????1????????????????????????????????????????????????????????????????:
        _15746_ = b[519:512];
      73'b???????1?????????????????????????????????????????????????????????????????:
        _15746_ = b[527:520];
      73'b??????1??????????????????????????????????????????????????????????????????:
        _15746_ = b[535:528];
      73'b?????1???????????????????????????????????????????????????????????????????:
        _15746_ = b[543:536];
      73'b????1????????????????????????????????????????????????????????????????????:
        _15746_ = b[551:544];
      73'b???1?????????????????????????????????????????????????????????????????????:
        _15746_ = b[559:552];
      73'b??1??????????????????????????????????????????????????????????????????????:
        _15746_ = b[567:560];
      73'b?1???????????????????????????????????????????????????????????????????????:
        _15746_ = b[575:568];
      73'b1????????????????????????????????????????????????????????????????????????:
        _15746_ = b[583:576];
      default:
        _15746_ = a;
    endcase
  endfunction
  assign vec_data_072 = _15746_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568], data_d1[583:576] }, { _06373_, _06372_, _06371_, _06370_, _06369_, _06368_, _06367_, _06366_, _06365_, _06364_, _06363_, _06362_, _06361_, _06360_, _06359_, _06358_, _06357_, _06356_, _06355_, _06354_, _06353_, _06352_, _06351_, _06350_, _06349_, _06348_, _06347_, _06346_, _06345_, _06344_, _06343_, _06342_, _06341_, _06340_, _06339_, _06338_, _06337_, _06336_, _06335_, _06334_, _06333_, _06332_, _06331_, _06330_, _06329_, _06328_, _06327_, _06326_, _06325_, _06324_, _06323_, _06322_, _06321_, _06320_, _06319_, _06318_, _06317_, _06316_, _06315_, _06314_, _06313_, _06312_, _06311_, _06310_, _06309_, _06308_, _06307_, _06306_, _06305_, _06304_, _06303_, _06302_, _06301_ });
  assign _06301_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1001001;
  assign _06302_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1001000;
  assign _06303_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000111;
  assign _06304_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000110;
  assign _06305_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000101;
  assign _06306_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000100;
  assign _06307_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000011;
  assign _06308_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000010;
  assign _06309_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000001;
  assign _06310_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 7'b1000000;
  assign _06311_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111111;
  assign _06312_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111110;
  assign _06313_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111101;
  assign _06314_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111100;
  assign _06315_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111011;
  assign _06316_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111010;
  assign _06317_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111001;
  assign _06318_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b111000;
  assign _06319_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110111;
  assign _06320_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110110;
  assign _06321_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110101;
  assign _06322_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110100;
  assign _06323_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110011;
  assign _06324_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110010;
  assign _06325_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110001;
  assign _06326_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b110000;
  assign _06327_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101111;
  assign _06328_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101110;
  assign _06329_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101101;
  assign _06330_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101100;
  assign _06331_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101011;
  assign _06332_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101010;
  assign _06333_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101001;
  assign _06334_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b101000;
  assign _06335_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100111;
  assign _06336_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100110;
  assign _06337_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100101;
  assign _06338_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100100;
  assign _06339_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7130|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100011;
  assign _06340_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7129|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100010;
  assign _06341_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7128|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100001;
  assign _06342_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7127|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 6'b100000;
  assign _06343_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7126|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11111;
  assign _06344_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11110;
  assign _06345_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11101;
  assign _06346_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11100;
  assign _06347_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11011;
  assign _06348_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11010;
  assign _06349_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11001;
  assign _06350_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b11000;
  assign _06351_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10111;
  assign _06352_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10110;
  assign _06353_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10101;
  assign _06354_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10100;
  assign _06355_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10011;
  assign _06356_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10010;
  assign _06357_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10001;
  assign _06358_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 5'b10000;
  assign _06359_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1111;
  assign _06360_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1110;
  assign _06361_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1101;
  assign _06362_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1100;
  assign _06363_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1011;
  assign _06364_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1010;
  assign _06365_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1001;
  assign _06366_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 4'b1000;
  assign _06367_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 3'b111;
  assign _06368_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 3'b110;
  assign _06369_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 3'b101;
  assign _06370_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 3'b100;
  assign _06371_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 2'b11;
  assign _06372_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 2'b10;
  assign _06373_ = vec_sum_072_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7095" *) 1'b1;
  function [7:0] _15820_;
    input [7:0] a;
    input [575:0] b;
    input [71:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *)
    (* parallel_case *)
    casez (s)
      72'b???????????????????????????????????????????????????????????????????????1:
        _15820_ = b[7:0];
      72'b??????????????????????????????????????????????????????????????????????1?:
        _15820_ = b[15:8];
      72'b?????????????????????????????????????????????????????????????????????1??:
        _15820_ = b[23:16];
      72'b????????????????????????????????????????????????????????????????????1???:
        _15820_ = b[31:24];
      72'b???????????????????????????????????????????????????????????????????1????:
        _15820_ = b[39:32];
      72'b??????????????????????????????????????????????????????????????????1?????:
        _15820_ = b[47:40];
      72'b?????????????????????????????????????????????????????????????????1??????:
        _15820_ = b[55:48];
      72'b????????????????????????????????????????????????????????????????1???????:
        _15820_ = b[63:56];
      72'b???????????????????????????????????????????????????????????????1????????:
        _15820_ = b[71:64];
      72'b??????????????????????????????????????????????????????????????1?????????:
        _15820_ = b[79:72];
      72'b?????????????????????????????????????????????????????????????1??????????:
        _15820_ = b[87:80];
      72'b????????????????????????????????????????????????????????????1???????????:
        _15820_ = b[95:88];
      72'b???????????????????????????????????????????????????????????1????????????:
        _15820_ = b[103:96];
      72'b??????????????????????????????????????????????????????????1?????????????:
        _15820_ = b[111:104];
      72'b?????????????????????????????????????????????????????????1??????????????:
        _15820_ = b[119:112];
      72'b????????????????????????????????????????????????????????1???????????????:
        _15820_ = b[127:120];
      72'b???????????????????????????????????????????????????????1????????????????:
        _15820_ = b[135:128];
      72'b??????????????????????????????????????????????????????1?????????????????:
        _15820_ = b[143:136];
      72'b?????????????????????????????????????????????????????1??????????????????:
        _15820_ = b[151:144];
      72'b????????????????????????????????????????????????????1???????????????????:
        _15820_ = b[159:152];
      72'b???????????????????????????????????????????????????1????????????????????:
        _15820_ = b[167:160];
      72'b??????????????????????????????????????????????????1?????????????????????:
        _15820_ = b[175:168];
      72'b?????????????????????????????????????????????????1??????????????????????:
        _15820_ = b[183:176];
      72'b????????????????????????????????????????????????1???????????????????????:
        _15820_ = b[191:184];
      72'b???????????????????????????????????????????????1????????????????????????:
        _15820_ = b[199:192];
      72'b??????????????????????????????????????????????1?????????????????????????:
        _15820_ = b[207:200];
      72'b?????????????????????????????????????????????1??????????????????????????:
        _15820_ = b[215:208];
      72'b????????????????????????????????????????????1???????????????????????????:
        _15820_ = b[223:216];
      72'b???????????????????????????????????????????1????????????????????????????:
        _15820_ = b[231:224];
      72'b??????????????????????????????????????????1?????????????????????????????:
        _15820_ = b[239:232];
      72'b?????????????????????????????????????????1??????????????????????????????:
        _15820_ = b[247:240];
      72'b????????????????????????????????????????1???????????????????????????????:
        _15820_ = b[255:248];
      72'b???????????????????????????????????????1????????????????????????????????:
        _15820_ = b[263:256];
      72'b??????????????????????????????????????1?????????????????????????????????:
        _15820_ = b[271:264];
      72'b?????????????????????????????????????1??????????????????????????????????:
        _15820_ = b[279:272];
      72'b????????????????????????????????????1???????????????????????????????????:
        _15820_ = b[287:280];
      72'b???????????????????????????????????1????????????????????????????????????:
        _15820_ = b[295:288];
      72'b??????????????????????????????????1?????????????????????????????????????:
        _15820_ = b[303:296];
      72'b?????????????????????????????????1??????????????????????????????????????:
        _15820_ = b[311:304];
      72'b????????????????????????????????1???????????????????????????????????????:
        _15820_ = b[319:312];
      72'b???????????????????????????????1????????????????????????????????????????:
        _15820_ = b[327:320];
      72'b??????????????????????????????1?????????????????????????????????????????:
        _15820_ = b[335:328];
      72'b?????????????????????????????1??????????????????????????????????????????:
        _15820_ = b[343:336];
      72'b????????????????????????????1???????????????????????????????????????????:
        _15820_ = b[351:344];
      72'b???????????????????????????1????????????????????????????????????????????:
        _15820_ = b[359:352];
      72'b??????????????????????????1?????????????????????????????????????????????:
        _15820_ = b[367:360];
      72'b?????????????????????????1??????????????????????????????????????????????:
        _15820_ = b[375:368];
      72'b????????????????????????1???????????????????????????????????????????????:
        _15820_ = b[383:376];
      72'b???????????????????????1????????????????????????????????????????????????:
        _15820_ = b[391:384];
      72'b??????????????????????1?????????????????????????????????????????????????:
        _15820_ = b[399:392];
      72'b?????????????????????1??????????????????????????????????????????????????:
        _15820_ = b[407:400];
      72'b????????????????????1???????????????????????????????????????????????????:
        _15820_ = b[415:408];
      72'b???????????????????1????????????????????????????????????????????????????:
        _15820_ = b[423:416];
      72'b??????????????????1?????????????????????????????????????????????????????:
        _15820_ = b[431:424];
      72'b?????????????????1??????????????????????????????????????????????????????:
        _15820_ = b[439:432];
      72'b????????????????1???????????????????????????????????????????????????????:
        _15820_ = b[447:440];
      72'b???????????????1????????????????????????????????????????????????????????:
        _15820_ = b[455:448];
      72'b??????????????1?????????????????????????????????????????????????????????:
        _15820_ = b[463:456];
      72'b?????????????1??????????????????????????????????????????????????????????:
        _15820_ = b[471:464];
      72'b????????????1???????????????????????????????????????????????????????????:
        _15820_ = b[479:472];
      72'b???????????1????????????????????????????????????????????????????????????:
        _15820_ = b[487:480];
      72'b??????????1?????????????????????????????????????????????????????????????:
        _15820_ = b[495:488];
      72'b?????????1??????????????????????????????????????????????????????????????:
        _15820_ = b[503:496];
      72'b????????1???????????????????????????????????????????????????????????????:
        _15820_ = b[511:504];
      72'b???????1????????????????????????????????????????????????????????????????:
        _15820_ = b[519:512];
      72'b??????1?????????????????????????????????????????????????????????????????:
        _15820_ = b[527:520];
      72'b?????1??????????????????????????????????????????????????????????????????:
        _15820_ = b[535:528];
      72'b????1???????????????????????????????????????????????????????????????????:
        _15820_ = b[543:536];
      72'b???1????????????????????????????????????????????????????????????????????:
        _15820_ = b[551:544];
      72'b??1?????????????????????????????????????????????????????????????????????:
        _15820_ = b[559:552];
      72'b?1??????????????????????????????????????????????????????????????????????:
        _15820_ = b[567:560];
      72'b1???????????????????????????????????????????????????????????????????????:
        _15820_ = b[575:568];
      default:
        _15820_ = a;
    endcase
  endfunction
  assign vec_data_071 = _15820_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560], data_d1[575:568] }, { _06445_, _06444_, _06443_, _06442_, _06441_, _06440_, _06439_, _06438_, _06437_, _06436_, _06435_, _06434_, _06433_, _06432_, _06431_, _06430_, _06429_, _06428_, _06427_, _06426_, _06425_, _06424_, _06423_, _06422_, _06421_, _06420_, _06419_, _06418_, _06417_, _06416_, _06415_, _06414_, _06413_, _06412_, _06411_, _06410_, _06409_, _06408_, _06407_, _06406_, _06405_, _06404_, _06403_, _06402_, _06401_, _06400_, _06399_, _06398_, _06397_, _06396_, _06395_, _06394_, _06393_, _06392_, _06391_, _06390_, _06389_, _06388_, _06387_, _06386_, _06385_, _06384_, _06383_, _06382_, _06381_, _06380_, _06379_, _06378_, _06377_, _06376_, _06375_, _06374_ });
  assign _06374_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1001000;
  assign _06375_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000111;
  assign _06376_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000110;
  assign _06377_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000101;
  assign _06378_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000100;
  assign _06379_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000011;
  assign _06380_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000010;
  assign _06381_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000001;
  assign _06382_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 7'b1000000;
  assign _06383_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111111;
  assign _06384_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111110;
  assign _06385_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111101;
  assign _06386_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111100;
  assign _06387_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111011;
  assign _06388_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111010;
  assign _06389_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111001;
  assign _06390_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b111000;
  assign _06391_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110111;
  assign _06392_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110110;
  assign _06393_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110101;
  assign _06394_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110100;
  assign _06395_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110011;
  assign _06396_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110010;
  assign _06397_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110001;
  assign _06398_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b110000;
  assign _06399_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101111;
  assign _06400_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101110;
  assign _06401_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101101;
  assign _06402_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101100;
  assign _06403_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101011;
  assign _06404_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101010;
  assign _06405_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101001;
  assign _06406_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b101000;
  assign _06407_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100111;
  assign _06408_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100110;
  assign _06409_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100101;
  assign _06410_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100100;
  assign _06411_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100011;
  assign _06412_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100010;
  assign _06413_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100001;
  assign _06414_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 6'b100000;
  assign _06415_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11111;
  assign _06416_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11110;
  assign _06417_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11101;
  assign _06418_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11100;
  assign _06419_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11011;
  assign _06420_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11010;
  assign _06421_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11001;
  assign _06422_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b11000;
  assign _06423_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10111;
  assign _06424_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10110;
  assign _06425_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10101;
  assign _06426_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10100;
  assign _06427_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10011;
  assign _06428_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10010;
  assign _06429_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10001;
  assign _06430_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 5'b10000;
  assign _06431_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1111;
  assign _06432_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1110;
  assign _06433_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1101;
  assign _06434_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1100;
  assign _06435_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1011;
  assign _06436_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1010;
  assign _06437_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1001;
  assign _06438_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 4'b1000;
  assign _06439_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 3'b111;
  assign _06440_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 3'b110;
  assign _06441_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 3'b101;
  assign _06442_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 3'b100;
  assign _06443_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 2'b11;
  assign _06444_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 2'b10;
  assign _06445_ = vec_sum_071_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7015" *) 1'b1;
  function [7:0] _15893_;
    input [7:0] a;
    input [567:0] b;
    input [70:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *)
    (* parallel_case *)
    casez (s)
      71'b??????????????????????????????????????????????????????????????????????1:
        _15893_ = b[7:0];
      71'b?????????????????????????????????????????????????????????????????????1?:
        _15893_ = b[15:8];
      71'b????????????????????????????????????????????????????????????????????1??:
        _15893_ = b[23:16];
      71'b???????????????????????????????????????????????????????????????????1???:
        _15893_ = b[31:24];
      71'b??????????????????????????????????????????????????????????????????1????:
        _15893_ = b[39:32];
      71'b?????????????????????????????????????????????????????????????????1?????:
        _15893_ = b[47:40];
      71'b????????????????????????????????????????????????????????????????1??????:
        _15893_ = b[55:48];
      71'b???????????????????????????????????????????????????????????????1???????:
        _15893_ = b[63:56];
      71'b??????????????????????????????????????????????????????????????1????????:
        _15893_ = b[71:64];
      71'b?????????????????????????????????????????????????????????????1?????????:
        _15893_ = b[79:72];
      71'b????????????????????????????????????????????????????????????1??????????:
        _15893_ = b[87:80];
      71'b???????????????????????????????????????????????????????????1???????????:
        _15893_ = b[95:88];
      71'b??????????????????????????????????????????????????????????1????????????:
        _15893_ = b[103:96];
      71'b?????????????????????????????????????????????????????????1?????????????:
        _15893_ = b[111:104];
      71'b????????????????????????????????????????????????????????1??????????????:
        _15893_ = b[119:112];
      71'b???????????????????????????????????????????????????????1???????????????:
        _15893_ = b[127:120];
      71'b??????????????????????????????????????????????????????1????????????????:
        _15893_ = b[135:128];
      71'b?????????????????????????????????????????????????????1?????????????????:
        _15893_ = b[143:136];
      71'b????????????????????????????????????????????????????1??????????????????:
        _15893_ = b[151:144];
      71'b???????????????????????????????????????????????????1???????????????????:
        _15893_ = b[159:152];
      71'b??????????????????????????????????????????????????1????????????????????:
        _15893_ = b[167:160];
      71'b?????????????????????????????????????????????????1?????????????????????:
        _15893_ = b[175:168];
      71'b????????????????????????????????????????????????1??????????????????????:
        _15893_ = b[183:176];
      71'b???????????????????????????????????????????????1???????????????????????:
        _15893_ = b[191:184];
      71'b??????????????????????????????????????????????1????????????????????????:
        _15893_ = b[199:192];
      71'b?????????????????????????????????????????????1?????????????????????????:
        _15893_ = b[207:200];
      71'b????????????????????????????????????????????1??????????????????????????:
        _15893_ = b[215:208];
      71'b???????????????????????????????????????????1???????????????????????????:
        _15893_ = b[223:216];
      71'b??????????????????????????????????????????1????????????????????????????:
        _15893_ = b[231:224];
      71'b?????????????????????????????????????????1?????????????????????????????:
        _15893_ = b[239:232];
      71'b????????????????????????????????????????1??????????????????????????????:
        _15893_ = b[247:240];
      71'b???????????????????????????????????????1???????????????????????????????:
        _15893_ = b[255:248];
      71'b??????????????????????????????????????1????????????????????????????????:
        _15893_ = b[263:256];
      71'b?????????????????????????????????????1?????????????????????????????????:
        _15893_ = b[271:264];
      71'b????????????????????????????????????1??????????????????????????????????:
        _15893_ = b[279:272];
      71'b???????????????????????????????????1???????????????????????????????????:
        _15893_ = b[287:280];
      71'b??????????????????????????????????1????????????????????????????????????:
        _15893_ = b[295:288];
      71'b?????????????????????????????????1?????????????????????????????????????:
        _15893_ = b[303:296];
      71'b????????????????????????????????1??????????????????????????????????????:
        _15893_ = b[311:304];
      71'b???????????????????????????????1???????????????????????????????????????:
        _15893_ = b[319:312];
      71'b??????????????????????????????1????????????????????????????????????????:
        _15893_ = b[327:320];
      71'b?????????????????????????????1?????????????????????????????????????????:
        _15893_ = b[335:328];
      71'b????????????????????????????1??????????????????????????????????????????:
        _15893_ = b[343:336];
      71'b???????????????????????????1???????????????????????????????????????????:
        _15893_ = b[351:344];
      71'b??????????????????????????1????????????????????????????????????????????:
        _15893_ = b[359:352];
      71'b?????????????????????????1?????????????????????????????????????????????:
        _15893_ = b[367:360];
      71'b????????????????????????1??????????????????????????????????????????????:
        _15893_ = b[375:368];
      71'b???????????????????????1???????????????????????????????????????????????:
        _15893_ = b[383:376];
      71'b??????????????????????1????????????????????????????????????????????????:
        _15893_ = b[391:384];
      71'b?????????????????????1?????????????????????????????????????????????????:
        _15893_ = b[399:392];
      71'b????????????????????1??????????????????????????????????????????????????:
        _15893_ = b[407:400];
      71'b???????????????????1???????????????????????????????????????????????????:
        _15893_ = b[415:408];
      71'b??????????????????1????????????????????????????????????????????????????:
        _15893_ = b[423:416];
      71'b?????????????????1?????????????????????????????????????????????????????:
        _15893_ = b[431:424];
      71'b????????????????1??????????????????????????????????????????????????????:
        _15893_ = b[439:432];
      71'b???????????????1???????????????????????????????????????????????????????:
        _15893_ = b[447:440];
      71'b??????????????1????????????????????????????????????????????????????????:
        _15893_ = b[455:448];
      71'b?????????????1?????????????????????????????????????????????????????????:
        _15893_ = b[463:456];
      71'b????????????1??????????????????????????????????????????????????????????:
        _15893_ = b[471:464];
      71'b???????????1???????????????????????????????????????????????????????????:
        _15893_ = b[479:472];
      71'b??????????1????????????????????????????????????????????????????????????:
        _15893_ = b[487:480];
      71'b?????????1?????????????????????????????????????????????????????????????:
        _15893_ = b[495:488];
      71'b????????1??????????????????????????????????????????????????????????????:
        _15893_ = b[503:496];
      71'b???????1???????????????????????????????????????????????????????????????:
        _15893_ = b[511:504];
      71'b??????1????????????????????????????????????????????????????????????????:
        _15893_ = b[519:512];
      71'b?????1?????????????????????????????????????????????????????????????????:
        _15893_ = b[527:520];
      71'b????1??????????????????????????????????????????????????????????????????:
        _15893_ = b[535:528];
      71'b???1???????????????????????????????????????????????????????????????????:
        _15893_ = b[543:536];
      71'b??1????????????????????????????????????????????????????????????????????:
        _15893_ = b[551:544];
      71'b?1?????????????????????????????????????????????????????????????????????:
        _15893_ = b[559:552];
      71'b1??????????????????????????????????????????????????????????????????????:
        _15893_ = b[567:560];
      default:
        _15893_ = a;
    endcase
  endfunction
  assign vec_data_070 = _15893_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552], data_d1[567:560] }, { _06516_, _06515_, _06514_, _06513_, _06512_, _06511_, _06510_, _06509_, _06508_, _06507_, _06506_, _06505_, _06504_, _06503_, _06502_, _06501_, _06500_, _06499_, _06498_, _06497_, _06496_, _06495_, _06494_, _06493_, _06492_, _06491_, _06490_, _06489_, _06488_, _06487_, _06486_, _06485_, _06484_, _06483_, _06482_, _06481_, _06480_, _06479_, _06478_, _06477_, _06476_, _06475_, _06474_, _06473_, _06472_, _06471_, _06470_, _06469_, _06468_, _06467_, _06466_, _06465_, _06464_, _06463_, _06462_, _06461_, _06460_, _06459_, _06458_, _06457_, _06456_, _06455_, _06454_, _06453_, _06452_, _06451_, _06450_, _06449_, _06448_, _06447_, _06446_ });
  assign _06446_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000111;
  assign _06447_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000110;
  assign _06448_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000101;
  assign _06449_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000100;
  assign _06450_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000011;
  assign _06451_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000010;
  assign _06452_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000001;
  assign _06453_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:7000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 7'b1000000;
  assign _06454_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111111;
  assign _06455_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111110;
  assign _06456_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111101;
  assign _06457_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111100;
  assign _06458_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111011;
  assign _06459_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111010;
  assign _06460_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111001;
  assign _06461_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b111000;
  assign _06462_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110111;
  assign _06463_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110110;
  assign _06464_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110101;
  assign _06465_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110100;
  assign _06466_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110011;
  assign _06467_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110010;
  assign _06468_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110001;
  assign _06469_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b110000;
  assign _06470_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101111;
  assign _06471_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101110;
  assign _06472_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101101;
  assign _06473_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101100;
  assign _06474_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101011;
  assign _06475_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101010;
  assign _06476_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101001;
  assign _06477_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b101000;
  assign _06478_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100111;
  assign _06479_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100110;
  assign _06480_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100101;
  assign _06481_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100100;
  assign _06482_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100011;
  assign _06483_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100010;
  assign _06484_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100001;
  assign _06485_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 6'b100000;
  assign _06486_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11111;
  assign _06487_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11110;
  assign _06488_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11101;
  assign _06489_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11100;
  assign _06490_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11011;
  assign _06491_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11010;
  assign _06492_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11001;
  assign _06493_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b11000;
  assign _06494_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10111;
  assign _06495_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10110;
  assign _06496_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10101;
  assign _06497_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10100;
  assign _06498_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10011;
  assign _06499_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10010;
  assign _06500_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10001;
  assign _06501_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 5'b10000;
  assign _06502_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1111;
  assign _06503_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1110;
  assign _06504_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1101;
  assign _06505_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1100;
  assign _06506_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1011;
  assign _06507_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1010;
  assign _06508_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1001;
  assign _06509_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 4'b1000;
  assign _06510_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 3'b111;
  assign _06511_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 3'b110;
  assign _06512_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 3'b101;
  assign _06513_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 3'b100;
  assign _06514_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 2'b11;
  assign _06515_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 2'b10;
  assign _06516_ = vec_sum_070_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6936" *) 1'b1;
  function [7:0] _15965_;
    input [7:0] a;
    input [559:0] b;
    input [69:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *)
    (* parallel_case *)
    casez (s)
      70'b?????????????????????????????????????????????????????????????????????1:
        _15965_ = b[7:0];
      70'b????????????????????????????????????????????????????????????????????1?:
        _15965_ = b[15:8];
      70'b???????????????????????????????????????????????????????????????????1??:
        _15965_ = b[23:16];
      70'b??????????????????????????????????????????????????????????????????1???:
        _15965_ = b[31:24];
      70'b?????????????????????????????????????????????????????????????????1????:
        _15965_ = b[39:32];
      70'b????????????????????????????????????????????????????????????????1?????:
        _15965_ = b[47:40];
      70'b???????????????????????????????????????????????????????????????1??????:
        _15965_ = b[55:48];
      70'b??????????????????????????????????????????????????????????????1???????:
        _15965_ = b[63:56];
      70'b?????????????????????????????????????????????????????????????1????????:
        _15965_ = b[71:64];
      70'b????????????????????????????????????????????????????????????1?????????:
        _15965_ = b[79:72];
      70'b???????????????????????????????????????????????????????????1??????????:
        _15965_ = b[87:80];
      70'b??????????????????????????????????????????????????????????1???????????:
        _15965_ = b[95:88];
      70'b?????????????????????????????????????????????????????????1????????????:
        _15965_ = b[103:96];
      70'b????????????????????????????????????????????????????????1?????????????:
        _15965_ = b[111:104];
      70'b???????????????????????????????????????????????????????1??????????????:
        _15965_ = b[119:112];
      70'b??????????????????????????????????????????????????????1???????????????:
        _15965_ = b[127:120];
      70'b?????????????????????????????????????????????????????1????????????????:
        _15965_ = b[135:128];
      70'b????????????????????????????????????????????????????1?????????????????:
        _15965_ = b[143:136];
      70'b???????????????????????????????????????????????????1??????????????????:
        _15965_ = b[151:144];
      70'b??????????????????????????????????????????????????1???????????????????:
        _15965_ = b[159:152];
      70'b?????????????????????????????????????????????????1????????????????????:
        _15965_ = b[167:160];
      70'b????????????????????????????????????????????????1?????????????????????:
        _15965_ = b[175:168];
      70'b???????????????????????????????????????????????1??????????????????????:
        _15965_ = b[183:176];
      70'b??????????????????????????????????????????????1???????????????????????:
        _15965_ = b[191:184];
      70'b?????????????????????????????????????????????1????????????????????????:
        _15965_ = b[199:192];
      70'b????????????????????????????????????????????1?????????????????????????:
        _15965_ = b[207:200];
      70'b???????????????????????????????????????????1??????????????????????????:
        _15965_ = b[215:208];
      70'b??????????????????????????????????????????1???????????????????????????:
        _15965_ = b[223:216];
      70'b?????????????????????????????????????????1????????????????????????????:
        _15965_ = b[231:224];
      70'b????????????????????????????????????????1?????????????????????????????:
        _15965_ = b[239:232];
      70'b???????????????????????????????????????1??????????????????????????????:
        _15965_ = b[247:240];
      70'b??????????????????????????????????????1???????????????????????????????:
        _15965_ = b[255:248];
      70'b?????????????????????????????????????1????????????????????????????????:
        _15965_ = b[263:256];
      70'b????????????????????????????????????1?????????????????????????????????:
        _15965_ = b[271:264];
      70'b???????????????????????????????????1??????????????????????????????????:
        _15965_ = b[279:272];
      70'b??????????????????????????????????1???????????????????????????????????:
        _15965_ = b[287:280];
      70'b?????????????????????????????????1????????????????????????????????????:
        _15965_ = b[295:288];
      70'b????????????????????????????????1?????????????????????????????????????:
        _15965_ = b[303:296];
      70'b???????????????????????????????1??????????????????????????????????????:
        _15965_ = b[311:304];
      70'b??????????????????????????????1???????????????????????????????????????:
        _15965_ = b[319:312];
      70'b?????????????????????????????1????????????????????????????????????????:
        _15965_ = b[327:320];
      70'b????????????????????????????1?????????????????????????????????????????:
        _15965_ = b[335:328];
      70'b???????????????????????????1??????????????????????????????????????????:
        _15965_ = b[343:336];
      70'b??????????????????????????1???????????????????????????????????????????:
        _15965_ = b[351:344];
      70'b?????????????????????????1????????????????????????????????????????????:
        _15965_ = b[359:352];
      70'b????????????????????????1?????????????????????????????????????????????:
        _15965_ = b[367:360];
      70'b???????????????????????1??????????????????????????????????????????????:
        _15965_ = b[375:368];
      70'b??????????????????????1???????????????????????????????????????????????:
        _15965_ = b[383:376];
      70'b?????????????????????1????????????????????????????????????????????????:
        _15965_ = b[391:384];
      70'b????????????????????1?????????????????????????????????????????????????:
        _15965_ = b[399:392];
      70'b???????????????????1??????????????????????????????????????????????????:
        _15965_ = b[407:400];
      70'b??????????????????1???????????????????????????????????????????????????:
        _15965_ = b[415:408];
      70'b?????????????????1????????????????????????????????????????????????????:
        _15965_ = b[423:416];
      70'b????????????????1?????????????????????????????????????????????????????:
        _15965_ = b[431:424];
      70'b???????????????1??????????????????????????????????????????????????????:
        _15965_ = b[439:432];
      70'b??????????????1???????????????????????????????????????????????????????:
        _15965_ = b[447:440];
      70'b?????????????1????????????????????????????????????????????????????????:
        _15965_ = b[455:448];
      70'b????????????1?????????????????????????????????????????????????????????:
        _15965_ = b[463:456];
      70'b???????????1??????????????????????????????????????????????????????????:
        _15965_ = b[471:464];
      70'b??????????1???????????????????????????????????????????????????????????:
        _15965_ = b[479:472];
      70'b?????????1????????????????????????????????????????????????????????????:
        _15965_ = b[487:480];
      70'b????????1?????????????????????????????????????????????????????????????:
        _15965_ = b[495:488];
      70'b???????1??????????????????????????????????????????????????????????????:
        _15965_ = b[503:496];
      70'b??????1???????????????????????????????????????????????????????????????:
        _15965_ = b[511:504];
      70'b?????1????????????????????????????????????????????????????????????????:
        _15965_ = b[519:512];
      70'b????1?????????????????????????????????????????????????????????????????:
        _15965_ = b[527:520];
      70'b???1??????????????????????????????????????????????????????????????????:
        _15965_ = b[535:528];
      70'b??1???????????????????????????????????????????????????????????????????:
        _15965_ = b[543:536];
      70'b?1????????????????????????????????????????????????????????????????????:
        _15965_ = b[551:544];
      70'b1?????????????????????????????????????????????????????????????????????:
        _15965_ = b[559:552];
      default:
        _15965_ = a;
    endcase
  endfunction
  assign vec_data_069 = _15965_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544], data_d1[559:552] }, { _06586_, _06585_, _06584_, _06583_, _06582_, _06581_, _06580_, _06579_, _06578_, _06577_, _06576_, _06575_, _06574_, _06573_, _06572_, _06571_, _06570_, _06569_, _06568_, _06567_, _06566_, _06565_, _06564_, _06563_, _06562_, _06561_, _06560_, _06559_, _06558_, _06557_, _06556_, _06555_, _06554_, _06553_, _06552_, _06551_, _06550_, _06549_, _06548_, _06547_, _06546_, _06545_, _06544_, _06543_, _06542_, _06541_, _06540_, _06539_, _06538_, _06537_, _06536_, _06535_, _06534_, _06533_, _06532_, _06531_, _06530_, _06529_, _06528_, _06527_, _06526_, _06525_, _06524_, _06523_, _06522_, _06521_, _06520_, _06519_, _06518_, _06517_ });
  assign _06517_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000110;
  assign _06518_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000101;
  assign _06519_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000100;
  assign _06520_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000011;
  assign _06521_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000010;
  assign _06522_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000001;
  assign _06523_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 7'b1000000;
  assign _06524_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111111;
  assign _06525_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111110;
  assign _06526_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111101;
  assign _06527_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111100;
  assign _06528_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111011;
  assign _06529_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111010;
  assign _06530_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111001;
  assign _06531_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b111000;
  assign _06532_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110111;
  assign _06533_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110110;
  assign _06534_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110101;
  assign _06535_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110100;
  assign _06536_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110011;
  assign _06537_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110010;
  assign _06538_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110001;
  assign _06539_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b110000;
  assign _06540_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101111;
  assign _06541_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101110;
  assign _06542_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101101;
  assign _06543_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101100;
  assign _06544_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101011;
  assign _06545_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101010;
  assign _06546_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101001;
  assign _06547_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b101000;
  assign _06548_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100111;
  assign _06549_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100110;
  assign _06550_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100101;
  assign _06551_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100100;
  assign _06552_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100011;
  assign _06553_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100010;
  assign _06554_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100001;
  assign _06555_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 6'b100000;
  assign _06556_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11111;
  assign _06557_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11110;
  assign _06558_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11101;
  assign _06559_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11100;
  assign _06560_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11011;
  assign _06561_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11010;
  assign _06562_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11001;
  assign _06563_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b11000;
  assign _06564_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10111;
  assign _06565_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10110;
  assign _06566_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10101;
  assign _06567_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10100;
  assign _06568_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10011;
  assign _06569_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10010;
  assign _06570_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10001;
  assign _06571_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 5'b10000;
  assign _06572_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1111;
  assign _06573_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1110;
  assign _06574_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1101;
  assign _06575_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1100;
  assign _06576_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1011;
  assign _06577_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1010;
  assign _06578_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1001;
  assign _06579_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 4'b1000;
  assign _06580_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 3'b111;
  assign _06581_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 3'b110;
  assign _06582_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 3'b101;
  assign _06583_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 3'b100;
  assign _06584_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 2'b11;
  assign _06585_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 2'b10;
  assign _06586_ = vec_sum_069_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6858" *) 1'b1;
  function [7:0] _16036_;
    input [7:0] a;
    input [551:0] b;
    input [68:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *)
    (* parallel_case *)
    casez (s)
      69'b????????????????????????????????????????????????????????????????????1:
        _16036_ = b[7:0];
      69'b???????????????????????????????????????????????????????????????????1?:
        _16036_ = b[15:8];
      69'b??????????????????????????????????????????????????????????????????1??:
        _16036_ = b[23:16];
      69'b?????????????????????????????????????????????????????????????????1???:
        _16036_ = b[31:24];
      69'b????????????????????????????????????????????????????????????????1????:
        _16036_ = b[39:32];
      69'b???????????????????????????????????????????????????????????????1?????:
        _16036_ = b[47:40];
      69'b??????????????????????????????????????????????????????????????1??????:
        _16036_ = b[55:48];
      69'b?????????????????????????????????????????????????????????????1???????:
        _16036_ = b[63:56];
      69'b????????????????????????????????????????????????????????????1????????:
        _16036_ = b[71:64];
      69'b???????????????????????????????????????????????????????????1?????????:
        _16036_ = b[79:72];
      69'b??????????????????????????????????????????????????????????1??????????:
        _16036_ = b[87:80];
      69'b?????????????????????????????????????????????????????????1???????????:
        _16036_ = b[95:88];
      69'b????????????????????????????????????????????????????????1????????????:
        _16036_ = b[103:96];
      69'b???????????????????????????????????????????????????????1?????????????:
        _16036_ = b[111:104];
      69'b??????????????????????????????????????????????????????1??????????????:
        _16036_ = b[119:112];
      69'b?????????????????????????????????????????????????????1???????????????:
        _16036_ = b[127:120];
      69'b????????????????????????????????????????????????????1????????????????:
        _16036_ = b[135:128];
      69'b???????????????????????????????????????????????????1?????????????????:
        _16036_ = b[143:136];
      69'b??????????????????????????????????????????????????1??????????????????:
        _16036_ = b[151:144];
      69'b?????????????????????????????????????????????????1???????????????????:
        _16036_ = b[159:152];
      69'b????????????????????????????????????????????????1????????????????????:
        _16036_ = b[167:160];
      69'b???????????????????????????????????????????????1?????????????????????:
        _16036_ = b[175:168];
      69'b??????????????????????????????????????????????1??????????????????????:
        _16036_ = b[183:176];
      69'b?????????????????????????????????????????????1???????????????????????:
        _16036_ = b[191:184];
      69'b????????????????????????????????????????????1????????????????????????:
        _16036_ = b[199:192];
      69'b???????????????????????????????????????????1?????????????????????????:
        _16036_ = b[207:200];
      69'b??????????????????????????????????????????1??????????????????????????:
        _16036_ = b[215:208];
      69'b?????????????????????????????????????????1???????????????????????????:
        _16036_ = b[223:216];
      69'b????????????????????????????????????????1????????????????????????????:
        _16036_ = b[231:224];
      69'b???????????????????????????????????????1?????????????????????????????:
        _16036_ = b[239:232];
      69'b??????????????????????????????????????1??????????????????????????????:
        _16036_ = b[247:240];
      69'b?????????????????????????????????????1???????????????????????????????:
        _16036_ = b[255:248];
      69'b????????????????????????????????????1????????????????????????????????:
        _16036_ = b[263:256];
      69'b???????????????????????????????????1?????????????????????????????????:
        _16036_ = b[271:264];
      69'b??????????????????????????????????1??????????????????????????????????:
        _16036_ = b[279:272];
      69'b?????????????????????????????????1???????????????????????????????????:
        _16036_ = b[287:280];
      69'b????????????????????????????????1????????????????????????????????????:
        _16036_ = b[295:288];
      69'b???????????????????????????????1?????????????????????????????????????:
        _16036_ = b[303:296];
      69'b??????????????????????????????1??????????????????????????????????????:
        _16036_ = b[311:304];
      69'b?????????????????????????????1???????????????????????????????????????:
        _16036_ = b[319:312];
      69'b????????????????????????????1????????????????????????????????????????:
        _16036_ = b[327:320];
      69'b???????????????????????????1?????????????????????????????????????????:
        _16036_ = b[335:328];
      69'b??????????????????????????1??????????????????????????????????????????:
        _16036_ = b[343:336];
      69'b?????????????????????????1???????????????????????????????????????????:
        _16036_ = b[351:344];
      69'b????????????????????????1????????????????????????????????????????????:
        _16036_ = b[359:352];
      69'b???????????????????????1?????????????????????????????????????????????:
        _16036_ = b[367:360];
      69'b??????????????????????1??????????????????????????????????????????????:
        _16036_ = b[375:368];
      69'b?????????????????????1???????????????????????????????????????????????:
        _16036_ = b[383:376];
      69'b????????????????????1????????????????????????????????????????????????:
        _16036_ = b[391:384];
      69'b???????????????????1?????????????????????????????????????????????????:
        _16036_ = b[399:392];
      69'b??????????????????1??????????????????????????????????????????????????:
        _16036_ = b[407:400];
      69'b?????????????????1???????????????????????????????????????????????????:
        _16036_ = b[415:408];
      69'b????????????????1????????????????????????????????????????????????????:
        _16036_ = b[423:416];
      69'b???????????????1?????????????????????????????????????????????????????:
        _16036_ = b[431:424];
      69'b??????????????1??????????????????????????????????????????????????????:
        _16036_ = b[439:432];
      69'b?????????????1???????????????????????????????????????????????????????:
        _16036_ = b[447:440];
      69'b????????????1????????????????????????????????????????????????????????:
        _16036_ = b[455:448];
      69'b???????????1?????????????????????????????????????????????????????????:
        _16036_ = b[463:456];
      69'b??????????1??????????????????????????????????????????????????????????:
        _16036_ = b[471:464];
      69'b?????????1???????????????????????????????????????????????????????????:
        _16036_ = b[479:472];
      69'b????????1????????????????????????????????????????????????????????????:
        _16036_ = b[487:480];
      69'b???????1?????????????????????????????????????????????????????????????:
        _16036_ = b[495:488];
      69'b??????1??????????????????????????????????????????????????????????????:
        _16036_ = b[503:496];
      69'b?????1???????????????????????????????????????????????????????????????:
        _16036_ = b[511:504];
      69'b????1????????????????????????????????????????????????????????????????:
        _16036_ = b[519:512];
      69'b???1?????????????????????????????????????????????????????????????????:
        _16036_ = b[527:520];
      69'b??1??????????????????????????????????????????????????????????????????:
        _16036_ = b[535:528];
      69'b?1???????????????????????????????????????????????????????????????????:
        _16036_ = b[543:536];
      69'b1????????????????????????????????????????????????????????????????????:
        _16036_ = b[551:544];
      default:
        _16036_ = a;
    endcase
  endfunction
  assign vec_data_068 = _16036_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536], data_d1[551:544] }, { _06655_, _06654_, _06653_, _06652_, _06651_, _06650_, _06649_, _06648_, _06647_, _06646_, _06645_, _06644_, _06643_, _06642_, _06641_, _06640_, _06639_, _06638_, _06637_, _06636_, _06635_, _06634_, _06633_, _06632_, _06631_, _06630_, _06629_, _06628_, _06627_, _06626_, _06625_, _06624_, _06623_, _06622_, _06621_, _06620_, _06619_, _06618_, _06617_, _06616_, _06615_, _06614_, _06613_, _06612_, _06611_, _06610_, _06609_, _06608_, _06607_, _06606_, _06605_, _06604_, _06603_, _06602_, _06601_, _06600_, _06599_, _06598_, _06597_, _06596_, _06595_, _06594_, _06593_, _06592_, _06591_, _06590_, _06589_, _06588_, _06587_ });
  assign _06587_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000101;
  assign _06588_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000100;
  assign _06589_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000011;
  assign _06590_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000010;
  assign _06591_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000001;
  assign _06592_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 7'b1000000;
  assign _06593_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111111;
  assign _06594_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111110;
  assign _06595_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111101;
  assign _06596_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111100;
  assign _06597_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111011;
  assign _06598_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111010;
  assign _06599_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111001;
  assign _06600_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b111000;
  assign _06601_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110111;
  assign _06602_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110110;
  assign _06603_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110101;
  assign _06604_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110100;
  assign _06605_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110011;
  assign _06606_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110010;
  assign _06607_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110001;
  assign _06608_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b110000;
  assign _06609_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101111;
  assign _06610_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101110;
  assign _06611_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101101;
  assign _06612_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101100;
  assign _06613_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101011;
  assign _06614_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101010;
  assign _06615_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101001;
  assign _06616_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b101000;
  assign _06617_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100111;
  assign _06618_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100110;
  assign _06619_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100101;
  assign _06620_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100100;
  assign _06621_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100011;
  assign _06622_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100010;
  assign _06623_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100001;
  assign _06624_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 6'b100000;
  assign _06625_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11111;
  assign _06626_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11110;
  assign _06627_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11101;
  assign _06628_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11100;
  assign _06629_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11011;
  assign _06630_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11010;
  assign _06631_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11001;
  assign _06632_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b11000;
  assign _06633_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10111;
  assign _06634_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10110;
  assign _06635_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10101;
  assign _06636_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6801|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10100;
  assign _06637_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10011;
  assign _06638_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10010;
  assign _06639_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10001;
  assign _06640_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 5'b10000;
  assign _06641_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1111;
  assign _06642_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1110;
  assign _06643_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1101;
  assign _06644_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1100;
  assign _06645_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1011;
  assign _06646_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1010;
  assign _06647_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1001;
  assign _06648_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 4'b1000;
  assign _06649_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 3'b111;
  assign _06650_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 3'b110;
  assign _06651_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 3'b101;
  assign _06652_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 3'b100;
  assign _06653_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 2'b11;
  assign _06654_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 2'b10;
  assign _06655_ = vec_sum_068_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6781" *) 1'b1;
  function [7:0] _16106_;
    input [7:0] a;
    input [543:0] b;
    input [67:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *)
    (* parallel_case *)
    casez (s)
      68'b???????????????????????????????????????????????????????????????????1:
        _16106_ = b[7:0];
      68'b??????????????????????????????????????????????????????????????????1?:
        _16106_ = b[15:8];
      68'b?????????????????????????????????????????????????????????????????1??:
        _16106_ = b[23:16];
      68'b????????????????????????????????????????????????????????????????1???:
        _16106_ = b[31:24];
      68'b???????????????????????????????????????????????????????????????1????:
        _16106_ = b[39:32];
      68'b??????????????????????????????????????????????????????????????1?????:
        _16106_ = b[47:40];
      68'b?????????????????????????????????????????????????????????????1??????:
        _16106_ = b[55:48];
      68'b????????????????????????????????????????????????????????????1???????:
        _16106_ = b[63:56];
      68'b???????????????????????????????????????????????????????????1????????:
        _16106_ = b[71:64];
      68'b??????????????????????????????????????????????????????????1?????????:
        _16106_ = b[79:72];
      68'b?????????????????????????????????????????????????????????1??????????:
        _16106_ = b[87:80];
      68'b????????????????????????????????????????????????????????1???????????:
        _16106_ = b[95:88];
      68'b???????????????????????????????????????????????????????1????????????:
        _16106_ = b[103:96];
      68'b??????????????????????????????????????????????????????1?????????????:
        _16106_ = b[111:104];
      68'b?????????????????????????????????????????????????????1??????????????:
        _16106_ = b[119:112];
      68'b????????????????????????????????????????????????????1???????????????:
        _16106_ = b[127:120];
      68'b???????????????????????????????????????????????????1????????????????:
        _16106_ = b[135:128];
      68'b??????????????????????????????????????????????????1?????????????????:
        _16106_ = b[143:136];
      68'b?????????????????????????????????????????????????1??????????????????:
        _16106_ = b[151:144];
      68'b????????????????????????????????????????????????1???????????????????:
        _16106_ = b[159:152];
      68'b???????????????????????????????????????????????1????????????????????:
        _16106_ = b[167:160];
      68'b??????????????????????????????????????????????1?????????????????????:
        _16106_ = b[175:168];
      68'b?????????????????????????????????????????????1??????????????????????:
        _16106_ = b[183:176];
      68'b????????????????????????????????????????????1???????????????????????:
        _16106_ = b[191:184];
      68'b???????????????????????????????????????????1????????????????????????:
        _16106_ = b[199:192];
      68'b??????????????????????????????????????????1?????????????????????????:
        _16106_ = b[207:200];
      68'b?????????????????????????????????????????1??????????????????????????:
        _16106_ = b[215:208];
      68'b????????????????????????????????????????1???????????????????????????:
        _16106_ = b[223:216];
      68'b???????????????????????????????????????1????????????????????????????:
        _16106_ = b[231:224];
      68'b??????????????????????????????????????1?????????????????????????????:
        _16106_ = b[239:232];
      68'b?????????????????????????????????????1??????????????????????????????:
        _16106_ = b[247:240];
      68'b????????????????????????????????????1???????????????????????????????:
        _16106_ = b[255:248];
      68'b???????????????????????????????????1????????????????????????????????:
        _16106_ = b[263:256];
      68'b??????????????????????????????????1?????????????????????????????????:
        _16106_ = b[271:264];
      68'b?????????????????????????????????1??????????????????????????????????:
        _16106_ = b[279:272];
      68'b????????????????????????????????1???????????????????????????????????:
        _16106_ = b[287:280];
      68'b???????????????????????????????1????????????????????????????????????:
        _16106_ = b[295:288];
      68'b??????????????????????????????1?????????????????????????????????????:
        _16106_ = b[303:296];
      68'b?????????????????????????????1??????????????????????????????????????:
        _16106_ = b[311:304];
      68'b????????????????????????????1???????????????????????????????????????:
        _16106_ = b[319:312];
      68'b???????????????????????????1????????????????????????????????????????:
        _16106_ = b[327:320];
      68'b??????????????????????????1?????????????????????????????????????????:
        _16106_ = b[335:328];
      68'b?????????????????????????1??????????????????????????????????????????:
        _16106_ = b[343:336];
      68'b????????????????????????1???????????????????????????????????????????:
        _16106_ = b[351:344];
      68'b???????????????????????1????????????????????????????????????????????:
        _16106_ = b[359:352];
      68'b??????????????????????1?????????????????????????????????????????????:
        _16106_ = b[367:360];
      68'b?????????????????????1??????????????????????????????????????????????:
        _16106_ = b[375:368];
      68'b????????????????????1???????????????????????????????????????????????:
        _16106_ = b[383:376];
      68'b???????????????????1????????????????????????????????????????????????:
        _16106_ = b[391:384];
      68'b??????????????????1?????????????????????????????????????????????????:
        _16106_ = b[399:392];
      68'b?????????????????1??????????????????????????????????????????????????:
        _16106_ = b[407:400];
      68'b????????????????1???????????????????????????????????????????????????:
        _16106_ = b[415:408];
      68'b???????????????1????????????????????????????????????????????????????:
        _16106_ = b[423:416];
      68'b??????????????1?????????????????????????????????????????????????????:
        _16106_ = b[431:424];
      68'b?????????????1??????????????????????????????????????????????????????:
        _16106_ = b[439:432];
      68'b????????????1???????????????????????????????????????????????????????:
        _16106_ = b[447:440];
      68'b???????????1????????????????????????????????????????????????????????:
        _16106_ = b[455:448];
      68'b??????????1?????????????????????????????????????????????????????????:
        _16106_ = b[463:456];
      68'b?????????1??????????????????????????????????????????????????????????:
        _16106_ = b[471:464];
      68'b????????1???????????????????????????????????????????????????????????:
        _16106_ = b[479:472];
      68'b???????1????????????????????????????????????????????????????????????:
        _16106_ = b[487:480];
      68'b??????1?????????????????????????????????????????????????????????????:
        _16106_ = b[495:488];
      68'b?????1??????????????????????????????????????????????????????????????:
        _16106_ = b[503:496];
      68'b????1???????????????????????????????????????????????????????????????:
        _16106_ = b[511:504];
      68'b???1????????????????????????????????????????????????????????????????:
        _16106_ = b[519:512];
      68'b??1?????????????????????????????????????????????????????????????????:
        _16106_ = b[527:520];
      68'b?1??????????????????????????????????????????????????????????????????:
        _16106_ = b[535:528];
      68'b1???????????????????????????????????????????????????????????????????:
        _16106_ = b[543:536];
      default:
        _16106_ = a;
    endcase
  endfunction
  assign vec_data_067 = _16106_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528], data_d1[543:536] }, { _06723_, _06722_, _06721_, _06720_, _06719_, _06718_, _06717_, _06716_, _06715_, _06714_, _06713_, _06712_, _06711_, _06710_, _06709_, _06708_, _06707_, _06706_, _06705_, _06704_, _06703_, _06702_, _06701_, _06700_, _06699_, _06698_, _06697_, _06696_, _06695_, _06694_, _06693_, _06692_, _06691_, _06690_, _06689_, _06688_, _06687_, _06686_, _06685_, _06684_, _06683_, _06682_, _06681_, _06680_, _06679_, _06678_, _06677_, _06676_, _06675_, _06674_, _06673_, _06672_, _06671_, _06670_, _06669_, _06668_, _06667_, _06666_, _06665_, _06664_, _06663_, _06662_, _06661_, _06660_, _06659_, _06658_, _06657_, _06656_ });
  assign _06656_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 7'b1000100;
  assign _06657_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 7'b1000011;
  assign _06658_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 7'b1000010;
  assign _06659_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 7'b1000001;
  assign _06660_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 7'b1000000;
  assign _06661_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111111;
  assign _06662_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111110;
  assign _06663_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111101;
  assign _06664_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111100;
  assign _06665_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111011;
  assign _06666_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111010;
  assign _06667_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111001;
  assign _06668_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b111000;
  assign _06669_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110111;
  assign _06670_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110110;
  assign _06671_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110101;
  assign _06672_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110100;
  assign _06673_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110011;
  assign _06674_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110010;
  assign _06675_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110001;
  assign _06676_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b110000;
  assign _06677_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101111;
  assign _06678_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101110;
  assign _06679_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101101;
  assign _06680_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101100;
  assign _06681_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101011;
  assign _06682_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101010;
  assign _06683_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101001;
  assign _06684_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b101000;
  assign _06685_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100111;
  assign _06686_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100110;
  assign _06687_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100101;
  assign _06688_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100100;
  assign _06689_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100011;
  assign _06690_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100010;
  assign _06691_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100001;
  assign _06692_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 6'b100000;
  assign _06693_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11111;
  assign _06694_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11110;
  assign _06695_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11101;
  assign _06696_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11100;
  assign _06697_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11011;
  assign _06698_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11010;
  assign _06699_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11001;
  assign _06700_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b11000;
  assign _06701_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10111;
  assign _06702_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10110;
  assign _06703_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10101;
  assign _06704_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10100;
  assign _06705_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10011;
  assign _06706_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10010;
  assign _06707_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10001;
  assign _06708_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 5'b10000;
  assign _06709_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1111;
  assign _06710_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1110;
  assign _06711_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1101;
  assign _06712_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1100;
  assign _06713_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1011;
  assign _06714_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1010;
  assign _06715_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1001;
  assign _06716_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 4'b1000;
  assign _06717_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 3'b111;
  assign _06718_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 3'b110;
  assign _06719_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 3'b101;
  assign _06720_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 3'b100;
  assign _06721_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 2'b11;
  assign _06722_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 2'b10;
  assign _06723_ = vec_sum_067_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6705" *) 1'b1;
  function [7:0] _16175_;
    input [7:0] a;
    input [535:0] b;
    input [66:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *)
    (* parallel_case *)
    casez (s)
      67'b??????????????????????????????????????????????????????????????????1:
        _16175_ = b[7:0];
      67'b?????????????????????????????????????????????????????????????????1?:
        _16175_ = b[15:8];
      67'b????????????????????????????????????????????????????????????????1??:
        _16175_ = b[23:16];
      67'b???????????????????????????????????????????????????????????????1???:
        _16175_ = b[31:24];
      67'b??????????????????????????????????????????????????????????????1????:
        _16175_ = b[39:32];
      67'b?????????????????????????????????????????????????????????????1?????:
        _16175_ = b[47:40];
      67'b????????????????????????????????????????????????????????????1??????:
        _16175_ = b[55:48];
      67'b???????????????????????????????????????????????????????????1???????:
        _16175_ = b[63:56];
      67'b??????????????????????????????????????????????????????????1????????:
        _16175_ = b[71:64];
      67'b?????????????????????????????????????????????????????????1?????????:
        _16175_ = b[79:72];
      67'b????????????????????????????????????????????????????????1??????????:
        _16175_ = b[87:80];
      67'b???????????????????????????????????????????????????????1???????????:
        _16175_ = b[95:88];
      67'b??????????????????????????????????????????????????????1????????????:
        _16175_ = b[103:96];
      67'b?????????????????????????????????????????????????????1?????????????:
        _16175_ = b[111:104];
      67'b????????????????????????????????????????????????????1??????????????:
        _16175_ = b[119:112];
      67'b???????????????????????????????????????????????????1???????????????:
        _16175_ = b[127:120];
      67'b??????????????????????????????????????????????????1????????????????:
        _16175_ = b[135:128];
      67'b?????????????????????????????????????????????????1?????????????????:
        _16175_ = b[143:136];
      67'b????????????????????????????????????????????????1??????????????????:
        _16175_ = b[151:144];
      67'b???????????????????????????????????????????????1???????????????????:
        _16175_ = b[159:152];
      67'b??????????????????????????????????????????????1????????????????????:
        _16175_ = b[167:160];
      67'b?????????????????????????????????????????????1?????????????????????:
        _16175_ = b[175:168];
      67'b????????????????????????????????????????????1??????????????????????:
        _16175_ = b[183:176];
      67'b???????????????????????????????????????????1???????????????????????:
        _16175_ = b[191:184];
      67'b??????????????????????????????????????????1????????????????????????:
        _16175_ = b[199:192];
      67'b?????????????????????????????????????????1?????????????????????????:
        _16175_ = b[207:200];
      67'b????????????????????????????????????????1??????????????????????????:
        _16175_ = b[215:208];
      67'b???????????????????????????????????????1???????????????????????????:
        _16175_ = b[223:216];
      67'b??????????????????????????????????????1????????????????????????????:
        _16175_ = b[231:224];
      67'b?????????????????????????????????????1?????????????????????????????:
        _16175_ = b[239:232];
      67'b????????????????????????????????????1??????????????????????????????:
        _16175_ = b[247:240];
      67'b???????????????????????????????????1???????????????????????????????:
        _16175_ = b[255:248];
      67'b??????????????????????????????????1????????????????????????????????:
        _16175_ = b[263:256];
      67'b?????????????????????????????????1?????????????????????????????????:
        _16175_ = b[271:264];
      67'b????????????????????????????????1??????????????????????????????????:
        _16175_ = b[279:272];
      67'b???????????????????????????????1???????????????????????????????????:
        _16175_ = b[287:280];
      67'b??????????????????????????????1????????????????????????????????????:
        _16175_ = b[295:288];
      67'b?????????????????????????????1?????????????????????????????????????:
        _16175_ = b[303:296];
      67'b????????????????????????????1??????????????????????????????????????:
        _16175_ = b[311:304];
      67'b???????????????????????????1???????????????????????????????????????:
        _16175_ = b[319:312];
      67'b??????????????????????????1????????????????????????????????????????:
        _16175_ = b[327:320];
      67'b?????????????????????????1?????????????????????????????????????????:
        _16175_ = b[335:328];
      67'b????????????????????????1??????????????????????????????????????????:
        _16175_ = b[343:336];
      67'b???????????????????????1???????????????????????????????????????????:
        _16175_ = b[351:344];
      67'b??????????????????????1????????????????????????????????????????????:
        _16175_ = b[359:352];
      67'b?????????????????????1?????????????????????????????????????????????:
        _16175_ = b[367:360];
      67'b????????????????????1??????????????????????????????????????????????:
        _16175_ = b[375:368];
      67'b???????????????????1???????????????????????????????????????????????:
        _16175_ = b[383:376];
      67'b??????????????????1????????????????????????????????????????????????:
        _16175_ = b[391:384];
      67'b?????????????????1?????????????????????????????????????????????????:
        _16175_ = b[399:392];
      67'b????????????????1??????????????????????????????????????????????????:
        _16175_ = b[407:400];
      67'b???????????????1???????????????????????????????????????????????????:
        _16175_ = b[415:408];
      67'b??????????????1????????????????????????????????????????????????????:
        _16175_ = b[423:416];
      67'b?????????????1?????????????????????????????????????????????????????:
        _16175_ = b[431:424];
      67'b????????????1??????????????????????????????????????????????????????:
        _16175_ = b[439:432];
      67'b???????????1???????????????????????????????????????????????????????:
        _16175_ = b[447:440];
      67'b??????????1????????????????????????????????????????????????????????:
        _16175_ = b[455:448];
      67'b?????????1?????????????????????????????????????????????????????????:
        _16175_ = b[463:456];
      67'b????????1??????????????????????????????????????????????????????????:
        _16175_ = b[471:464];
      67'b???????1???????????????????????????????????????????????????????????:
        _16175_ = b[479:472];
      67'b??????1????????????????????????????????????????????????????????????:
        _16175_ = b[487:480];
      67'b?????1?????????????????????????????????????????????????????????????:
        _16175_ = b[495:488];
      67'b????1??????????????????????????????????????????????????????????????:
        _16175_ = b[503:496];
      67'b???1???????????????????????????????????????????????????????????????:
        _16175_ = b[511:504];
      67'b??1????????????????????????????????????????????????????????????????:
        _16175_ = b[519:512];
      67'b?1?????????????????????????????????????????????????????????????????:
        _16175_ = b[527:520];
      67'b1??????????????????????????????????????????????????????????????????:
        _16175_ = b[535:528];
      default:
        _16175_ = a;
    endcase
  endfunction
  assign vec_data_066 = _16175_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520], data_d1[535:528] }, { _06790_, _06789_, _06788_, _06787_, _06786_, _06785_, _06784_, _06783_, _06782_, _06781_, _06780_, _06779_, _06778_, _06777_, _06776_, _06775_, _06774_, _06773_, _06772_, _06771_, _06770_, _06769_, _06768_, _06767_, _06766_, _06765_, _06764_, _06763_, _06762_, _06761_, _06760_, _06759_, _06758_, _06757_, _06756_, _06755_, _06754_, _06753_, _06752_, _06751_, _06750_, _06749_, _06748_, _06747_, _06746_, _06745_, _06744_, _06743_, _06742_, _06741_, _06740_, _06739_, _06738_, _06737_, _06736_, _06735_, _06734_, _06733_, _06732_, _06731_, _06730_, _06729_, _06728_, _06727_, _06726_, _06725_, _06724_ });
  assign _06724_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 7'b1000011;
  assign _06725_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 7'b1000010;
  assign _06726_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 7'b1000001;
  assign _06727_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 7'b1000000;
  assign _06728_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111111;
  assign _06729_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111110;
  assign _06730_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111101;
  assign _06731_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111100;
  assign _06732_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111011;
  assign _06733_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111010;
  assign _06734_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111001;
  assign _06735_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b111000;
  assign _06736_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110111;
  assign _06737_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110110;
  assign _06738_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110101;
  assign _06739_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110100;
  assign _06740_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110011;
  assign _06741_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110010;
  assign _06742_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110001;
  assign _06743_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b110000;
  assign _06744_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101111;
  assign _06745_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101110;
  assign _06746_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101101;
  assign _06747_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101100;
  assign _06748_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101011;
  assign _06749_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101010;
  assign _06750_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101001;
  assign _06751_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b101000;
  assign _06752_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100111;
  assign _06753_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100110;
  assign _06754_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100101;
  assign _06755_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100100;
  assign _06756_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100011;
  assign _06757_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100010;
  assign _06758_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100001;
  assign _06759_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 6'b100000;
  assign _06760_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11111;
  assign _06761_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11110;
  assign _06762_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11101;
  assign _06763_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11100;
  assign _06764_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11011;
  assign _06765_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11010;
  assign _06766_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11001;
  assign _06767_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b11000;
  assign _06768_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10111;
  assign _06769_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10110;
  assign _06770_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10101;
  assign _06771_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10100;
  assign _06772_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10011;
  assign _06773_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10010;
  assign _06774_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10001;
  assign _06775_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 5'b10000;
  assign _06776_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1111;
  assign _06777_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1110;
  assign _06778_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1101;
  assign _06779_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1100;
  assign _06780_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1011;
  assign _06781_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1010;
  assign _06782_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1001;
  assign _06783_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 4'b1000;
  assign _06784_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 3'b111;
  assign _06785_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 3'b110;
  assign _06786_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 3'b101;
  assign _06787_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 3'b100;
  assign _06788_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 2'b11;
  assign _06789_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 2'b10;
  assign _06790_ = vec_sum_066_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6630" *) 1'b1;
  function [7:0] _16243_;
    input [7:0] a;
    input [527:0] b;
    input [65:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *)
    (* parallel_case *)
    casez (s)
      66'b?????????????????????????????????????????????????????????????????1:
        _16243_ = b[7:0];
      66'b????????????????????????????????????????????????????????????????1?:
        _16243_ = b[15:8];
      66'b???????????????????????????????????????????????????????????????1??:
        _16243_ = b[23:16];
      66'b??????????????????????????????????????????????????????????????1???:
        _16243_ = b[31:24];
      66'b?????????????????????????????????????????????????????????????1????:
        _16243_ = b[39:32];
      66'b????????????????????????????????????????????????????????????1?????:
        _16243_ = b[47:40];
      66'b???????????????????????????????????????????????????????????1??????:
        _16243_ = b[55:48];
      66'b??????????????????????????????????????????????????????????1???????:
        _16243_ = b[63:56];
      66'b?????????????????????????????????????????????????????????1????????:
        _16243_ = b[71:64];
      66'b????????????????????????????????????????????????????????1?????????:
        _16243_ = b[79:72];
      66'b???????????????????????????????????????????????????????1??????????:
        _16243_ = b[87:80];
      66'b??????????????????????????????????????????????????????1???????????:
        _16243_ = b[95:88];
      66'b?????????????????????????????????????????????????????1????????????:
        _16243_ = b[103:96];
      66'b????????????????????????????????????????????????????1?????????????:
        _16243_ = b[111:104];
      66'b???????????????????????????????????????????????????1??????????????:
        _16243_ = b[119:112];
      66'b??????????????????????????????????????????????????1???????????????:
        _16243_ = b[127:120];
      66'b?????????????????????????????????????????????????1????????????????:
        _16243_ = b[135:128];
      66'b????????????????????????????????????????????????1?????????????????:
        _16243_ = b[143:136];
      66'b???????????????????????????????????????????????1??????????????????:
        _16243_ = b[151:144];
      66'b??????????????????????????????????????????????1???????????????????:
        _16243_ = b[159:152];
      66'b?????????????????????????????????????????????1????????????????????:
        _16243_ = b[167:160];
      66'b????????????????????????????????????????????1?????????????????????:
        _16243_ = b[175:168];
      66'b???????????????????????????????????????????1??????????????????????:
        _16243_ = b[183:176];
      66'b??????????????????????????????????????????1???????????????????????:
        _16243_ = b[191:184];
      66'b?????????????????????????????????????????1????????????????????????:
        _16243_ = b[199:192];
      66'b????????????????????????????????????????1?????????????????????????:
        _16243_ = b[207:200];
      66'b???????????????????????????????????????1??????????????????????????:
        _16243_ = b[215:208];
      66'b??????????????????????????????????????1???????????????????????????:
        _16243_ = b[223:216];
      66'b?????????????????????????????????????1????????????????????????????:
        _16243_ = b[231:224];
      66'b????????????????????????????????????1?????????????????????????????:
        _16243_ = b[239:232];
      66'b???????????????????????????????????1??????????????????????????????:
        _16243_ = b[247:240];
      66'b??????????????????????????????????1???????????????????????????????:
        _16243_ = b[255:248];
      66'b?????????????????????????????????1????????????????????????????????:
        _16243_ = b[263:256];
      66'b????????????????????????????????1?????????????????????????????????:
        _16243_ = b[271:264];
      66'b???????????????????????????????1??????????????????????????????????:
        _16243_ = b[279:272];
      66'b??????????????????????????????1???????????????????????????????????:
        _16243_ = b[287:280];
      66'b?????????????????????????????1????????????????????????????????????:
        _16243_ = b[295:288];
      66'b????????????????????????????1?????????????????????????????????????:
        _16243_ = b[303:296];
      66'b???????????????????????????1??????????????????????????????????????:
        _16243_ = b[311:304];
      66'b??????????????????????????1???????????????????????????????????????:
        _16243_ = b[319:312];
      66'b?????????????????????????1????????????????????????????????????????:
        _16243_ = b[327:320];
      66'b????????????????????????1?????????????????????????????????????????:
        _16243_ = b[335:328];
      66'b???????????????????????1??????????????????????????????????????????:
        _16243_ = b[343:336];
      66'b??????????????????????1???????????????????????????????????????????:
        _16243_ = b[351:344];
      66'b?????????????????????1????????????????????????????????????????????:
        _16243_ = b[359:352];
      66'b????????????????????1?????????????????????????????????????????????:
        _16243_ = b[367:360];
      66'b???????????????????1??????????????????????????????????????????????:
        _16243_ = b[375:368];
      66'b??????????????????1???????????????????????????????????????????????:
        _16243_ = b[383:376];
      66'b?????????????????1????????????????????????????????????????????????:
        _16243_ = b[391:384];
      66'b????????????????1?????????????????????????????????????????????????:
        _16243_ = b[399:392];
      66'b???????????????1??????????????????????????????????????????????????:
        _16243_ = b[407:400];
      66'b??????????????1???????????????????????????????????????????????????:
        _16243_ = b[415:408];
      66'b?????????????1????????????????????????????????????????????????????:
        _16243_ = b[423:416];
      66'b????????????1?????????????????????????????????????????????????????:
        _16243_ = b[431:424];
      66'b???????????1??????????????????????????????????????????????????????:
        _16243_ = b[439:432];
      66'b??????????1???????????????????????????????????????????????????????:
        _16243_ = b[447:440];
      66'b?????????1????????????????????????????????????????????????????????:
        _16243_ = b[455:448];
      66'b????????1?????????????????????????????????????????????????????????:
        _16243_ = b[463:456];
      66'b???????1??????????????????????????????????????????????????????????:
        _16243_ = b[471:464];
      66'b??????1???????????????????????????????????????????????????????????:
        _16243_ = b[479:472];
      66'b?????1????????????????????????????????????????????????????????????:
        _16243_ = b[487:480];
      66'b????1?????????????????????????????????????????????????????????????:
        _16243_ = b[495:488];
      66'b???1??????????????????????????????????????????????????????????????:
        _16243_ = b[503:496];
      66'b??1???????????????????????????????????????????????????????????????:
        _16243_ = b[511:504];
      66'b?1????????????????????????????????????????????????????????????????:
        _16243_ = b[519:512];
      66'b1?????????????????????????????????????????????????????????????????:
        _16243_ = b[527:520];
      default:
        _16243_ = a;
    endcase
  endfunction
  assign vec_data_065 = _16243_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512], data_d1[527:520] }, { _06856_, _06855_, _06854_, _06853_, _06852_, _06851_, _06850_, _06849_, _06848_, _06847_, _06846_, _06845_, _06844_, _06843_, _06842_, _06841_, _06840_, _06839_, _06838_, _06837_, _06836_, _06835_, _06834_, _06833_, _06832_, _06831_, _06830_, _06829_, _06828_, _06827_, _06826_, _06825_, _06824_, _06823_, _06822_, _06821_, _06820_, _06819_, _06818_, _06817_, _06816_, _06815_, _06814_, _06813_, _06812_, _06811_, _06810_, _06809_, _06808_, _06807_, _06806_, _06805_, _06804_, _06803_, _06802_, _06801_, _06800_, _06799_, _06798_, _06797_, _06796_, _06795_, _06794_, _06793_, _06792_, _06791_ });
  assign _06791_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 7'b1000010;
  assign _06792_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 7'b1000001;
  assign _06793_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 7'b1000000;
  assign _06794_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111111;
  assign _06795_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111110;
  assign _06796_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111101;
  assign _06797_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111100;
  assign _06798_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111011;
  assign _06799_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111010;
  assign _06800_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111001;
  assign _06801_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b111000;
  assign _06802_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110111;
  assign _06803_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110110;
  assign _06804_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110101;
  assign _06805_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110100;
  assign _06806_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110011;
  assign _06807_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110010;
  assign _06808_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110001;
  assign _06809_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b110000;
  assign _06810_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101111;
  assign _06811_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101110;
  assign _06812_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101101;
  assign _06813_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101100;
  assign _06814_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101011;
  assign _06815_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101010;
  assign _06816_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101001;
  assign _06817_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b101000;
  assign _06818_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100111;
  assign _06819_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100110;
  assign _06820_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100101;
  assign _06821_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100100;
  assign _06822_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100011;
  assign _06823_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100010;
  assign _06824_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100001;
  assign _06825_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 6'b100000;
  assign _06826_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11111;
  assign _06827_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11110;
  assign _06828_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11101;
  assign _06829_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11100;
  assign _06830_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11011;
  assign _06831_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11010;
  assign _06832_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11001;
  assign _06833_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b11000;
  assign _06834_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10111;
  assign _06835_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10110;
  assign _06836_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10101;
  assign _06837_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10100;
  assign _06838_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10011;
  assign _06839_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10010;
  assign _06840_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10001;
  assign _06841_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 5'b10000;
  assign _06842_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1111;
  assign _06843_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1110;
  assign _06844_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1101;
  assign _06845_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1100;
  assign _06846_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1011;
  assign _06847_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1010;
  assign _06848_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1001;
  assign _06849_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 4'b1000;
  assign _06850_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 3'b111;
  assign _06851_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 3'b110;
  assign _06852_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 3'b101;
  assign _06853_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 3'b100;
  assign _06854_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 2'b11;
  assign _06855_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 2'b10;
  assign _06856_ = vec_sum_065_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6556" *) 1'b1;
  function [7:0] _16310_;
    input [7:0] a;
    input [519:0] b;
    input [64:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *)
    (* parallel_case *)
    casez (s)
      65'b????????????????????????????????????????????????????????????????1:
        _16310_ = b[7:0];
      65'b???????????????????????????????????????????????????????????????1?:
        _16310_ = b[15:8];
      65'b??????????????????????????????????????????????????????????????1??:
        _16310_ = b[23:16];
      65'b?????????????????????????????????????????????????????????????1???:
        _16310_ = b[31:24];
      65'b????????????????????????????????????????????????????????????1????:
        _16310_ = b[39:32];
      65'b???????????????????????????????????????????????????????????1?????:
        _16310_ = b[47:40];
      65'b??????????????????????????????????????????????????????????1??????:
        _16310_ = b[55:48];
      65'b?????????????????????????????????????????????????????????1???????:
        _16310_ = b[63:56];
      65'b????????????????????????????????????????????????????????1????????:
        _16310_ = b[71:64];
      65'b???????????????????????????????????????????????????????1?????????:
        _16310_ = b[79:72];
      65'b??????????????????????????????????????????????????????1??????????:
        _16310_ = b[87:80];
      65'b?????????????????????????????????????????????????????1???????????:
        _16310_ = b[95:88];
      65'b????????????????????????????????????????????????????1????????????:
        _16310_ = b[103:96];
      65'b???????????????????????????????????????????????????1?????????????:
        _16310_ = b[111:104];
      65'b??????????????????????????????????????????????????1??????????????:
        _16310_ = b[119:112];
      65'b?????????????????????????????????????????????????1???????????????:
        _16310_ = b[127:120];
      65'b????????????????????????????????????????????????1????????????????:
        _16310_ = b[135:128];
      65'b???????????????????????????????????????????????1?????????????????:
        _16310_ = b[143:136];
      65'b??????????????????????????????????????????????1??????????????????:
        _16310_ = b[151:144];
      65'b?????????????????????????????????????????????1???????????????????:
        _16310_ = b[159:152];
      65'b????????????????????????????????????????????1????????????????????:
        _16310_ = b[167:160];
      65'b???????????????????????????????????????????1?????????????????????:
        _16310_ = b[175:168];
      65'b??????????????????????????????????????????1??????????????????????:
        _16310_ = b[183:176];
      65'b?????????????????????????????????????????1???????????????????????:
        _16310_ = b[191:184];
      65'b????????????????????????????????????????1????????????????????????:
        _16310_ = b[199:192];
      65'b???????????????????????????????????????1?????????????????????????:
        _16310_ = b[207:200];
      65'b??????????????????????????????????????1??????????????????????????:
        _16310_ = b[215:208];
      65'b?????????????????????????????????????1???????????????????????????:
        _16310_ = b[223:216];
      65'b????????????????????????????????????1????????????????????????????:
        _16310_ = b[231:224];
      65'b???????????????????????????????????1?????????????????????????????:
        _16310_ = b[239:232];
      65'b??????????????????????????????????1??????????????????????????????:
        _16310_ = b[247:240];
      65'b?????????????????????????????????1???????????????????????????????:
        _16310_ = b[255:248];
      65'b????????????????????????????????1????????????????????????????????:
        _16310_ = b[263:256];
      65'b???????????????????????????????1?????????????????????????????????:
        _16310_ = b[271:264];
      65'b??????????????????????????????1??????????????????????????????????:
        _16310_ = b[279:272];
      65'b?????????????????????????????1???????????????????????????????????:
        _16310_ = b[287:280];
      65'b????????????????????????????1????????????????????????????????????:
        _16310_ = b[295:288];
      65'b???????????????????????????1?????????????????????????????????????:
        _16310_ = b[303:296];
      65'b??????????????????????????1??????????????????????????????????????:
        _16310_ = b[311:304];
      65'b?????????????????????????1???????????????????????????????????????:
        _16310_ = b[319:312];
      65'b????????????????????????1????????????????????????????????????????:
        _16310_ = b[327:320];
      65'b???????????????????????1?????????????????????????????????????????:
        _16310_ = b[335:328];
      65'b??????????????????????1??????????????????????????????????????????:
        _16310_ = b[343:336];
      65'b?????????????????????1???????????????????????????????????????????:
        _16310_ = b[351:344];
      65'b????????????????????1????????????????????????????????????????????:
        _16310_ = b[359:352];
      65'b???????????????????1?????????????????????????????????????????????:
        _16310_ = b[367:360];
      65'b??????????????????1??????????????????????????????????????????????:
        _16310_ = b[375:368];
      65'b?????????????????1???????????????????????????????????????????????:
        _16310_ = b[383:376];
      65'b????????????????1????????????????????????????????????????????????:
        _16310_ = b[391:384];
      65'b???????????????1?????????????????????????????????????????????????:
        _16310_ = b[399:392];
      65'b??????????????1??????????????????????????????????????????????????:
        _16310_ = b[407:400];
      65'b?????????????1???????????????????????????????????????????????????:
        _16310_ = b[415:408];
      65'b????????????1????????????????????????????????????????????????????:
        _16310_ = b[423:416];
      65'b???????????1?????????????????????????????????????????????????????:
        _16310_ = b[431:424];
      65'b??????????1??????????????????????????????????????????????????????:
        _16310_ = b[439:432];
      65'b?????????1???????????????????????????????????????????????????????:
        _16310_ = b[447:440];
      65'b????????1????????????????????????????????????????????????????????:
        _16310_ = b[455:448];
      65'b???????1?????????????????????????????????????????????????????????:
        _16310_ = b[463:456];
      65'b??????1??????????????????????????????????????????????????????????:
        _16310_ = b[471:464];
      65'b?????1???????????????????????????????????????????????????????????:
        _16310_ = b[479:472];
      65'b????1????????????????????????????????????????????????????????????:
        _16310_ = b[487:480];
      65'b???1?????????????????????????????????????????????????????????????:
        _16310_ = b[495:488];
      65'b??1??????????????????????????????????????????????????????????????:
        _16310_ = b[503:496];
      65'b?1???????????????????????????????????????????????????????????????:
        _16310_ = b[511:504];
      65'b1????????????????????????????????????????????????????????????????:
        _16310_ = b[519:512];
      default:
        _16310_ = a;
    endcase
  endfunction
  assign vec_data_064 = _16310_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504], data_d1[519:512] }, { _06921_, _06920_, _06919_, _06918_, _06917_, _06916_, _06915_, _06914_, _06913_, _06912_, _06911_, _06910_, _06909_, _06908_, _06907_, _06906_, _06905_, _06904_, _06903_, _06902_, _06901_, _06900_, _06899_, _06898_, _06897_, _06896_, _06895_, _06894_, _06893_, _06892_, _06891_, _06890_, _06889_, _06888_, _06887_, _06886_, _06885_, _06884_, _06883_, _06882_, _06881_, _06880_, _06879_, _06878_, _06877_, _06876_, _06875_, _06874_, _06873_, _06872_, _06871_, _06870_, _06869_, _06868_, _06867_, _06866_, _06865_, _06864_, _06863_, _06862_, _06861_, _06860_, _06859_, _06858_, _06857_ });
  assign _06857_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 7'b1000001;
  assign _06858_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 7'b1000000;
  assign _06859_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111111;
  assign _06860_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111110;
  assign _06861_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111101;
  assign _06862_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111100;
  assign _06863_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111011;
  assign _06864_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111010;
  assign _06865_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111001;
  assign _06866_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b111000;
  assign _06867_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110111;
  assign _06868_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110110;
  assign _06869_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110101;
  assign _06870_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110100;
  assign _06871_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110011;
  assign _06872_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110010;
  assign _06873_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110001;
  assign _06874_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b110000;
  assign _06875_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101111;
  assign _06876_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101110;
  assign _06877_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101101;
  assign _06878_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101100;
  assign _06879_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101011;
  assign _06880_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101010;
  assign _06881_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101001;
  assign _06882_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b101000;
  assign _06883_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100111;
  assign _06884_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100110;
  assign _06885_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100101;
  assign _06886_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100100;
  assign _06887_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100011;
  assign _06888_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100010;
  assign _06889_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100001;
  assign _06890_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 6'b100000;
  assign _06891_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11111;
  assign _06892_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11110;
  assign _06893_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11101;
  assign _06894_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11100;
  assign _06895_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11011;
  assign _06896_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11010;
  assign _06897_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11001;
  assign _06898_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b11000;
  assign _06899_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10111;
  assign _06900_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10110;
  assign _06901_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10101;
  assign _06902_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10100;
  assign _06903_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10011;
  assign _06904_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10010;
  assign _06905_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10001;
  assign _06906_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 5'b10000;
  assign _06907_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1111;
  assign _06908_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1110;
  assign _06909_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1101;
  assign _06910_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1100;
  assign _06911_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1011;
  assign _06912_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1010;
  assign _06913_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1001;
  assign _06914_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 4'b1000;
  assign _06915_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 3'b111;
  assign _06916_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 3'b110;
  assign _06917_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 3'b101;
  assign _06918_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 3'b100;
  assign _06919_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 2'b11;
  assign _06920_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 2'b10;
  assign _06921_ = vec_sum_064_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6483" *) 1'b1;
  function [7:0] _16376_;
    input [7:0] a;
    input [511:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _16376_ = b[7:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _16376_ = b[15:8];
      64'b?????????????????????????????????????????????????????????????1??:
        _16376_ = b[23:16];
      64'b????????????????????????????????????????????????????????????1???:
        _16376_ = b[31:24];
      64'b???????????????????????????????????????????????????????????1????:
        _16376_ = b[39:32];
      64'b??????????????????????????????????????????????????????????1?????:
        _16376_ = b[47:40];
      64'b?????????????????????????????????????????????????????????1??????:
        _16376_ = b[55:48];
      64'b????????????????????????????????????????????????????????1???????:
        _16376_ = b[63:56];
      64'b???????????????????????????????????????????????????????1????????:
        _16376_ = b[71:64];
      64'b??????????????????????????????????????????????????????1?????????:
        _16376_ = b[79:72];
      64'b?????????????????????????????????????????????????????1??????????:
        _16376_ = b[87:80];
      64'b????????????????????????????????????????????????????1???????????:
        _16376_ = b[95:88];
      64'b???????????????????????????????????????????????????1????????????:
        _16376_ = b[103:96];
      64'b??????????????????????????????????????????????????1?????????????:
        _16376_ = b[111:104];
      64'b?????????????????????????????????????????????????1??????????????:
        _16376_ = b[119:112];
      64'b????????????????????????????????????????????????1???????????????:
        _16376_ = b[127:120];
      64'b???????????????????????????????????????????????1????????????????:
        _16376_ = b[135:128];
      64'b??????????????????????????????????????????????1?????????????????:
        _16376_ = b[143:136];
      64'b?????????????????????????????????????????????1??????????????????:
        _16376_ = b[151:144];
      64'b????????????????????????????????????????????1???????????????????:
        _16376_ = b[159:152];
      64'b???????????????????????????????????????????1????????????????????:
        _16376_ = b[167:160];
      64'b??????????????????????????????????????????1?????????????????????:
        _16376_ = b[175:168];
      64'b?????????????????????????????????????????1??????????????????????:
        _16376_ = b[183:176];
      64'b????????????????????????????????????????1???????????????????????:
        _16376_ = b[191:184];
      64'b???????????????????????????????????????1????????????????????????:
        _16376_ = b[199:192];
      64'b??????????????????????????????????????1?????????????????????????:
        _16376_ = b[207:200];
      64'b?????????????????????????????????????1??????????????????????????:
        _16376_ = b[215:208];
      64'b????????????????????????????????????1???????????????????????????:
        _16376_ = b[223:216];
      64'b???????????????????????????????????1????????????????????????????:
        _16376_ = b[231:224];
      64'b??????????????????????????????????1?????????????????????????????:
        _16376_ = b[239:232];
      64'b?????????????????????????????????1??????????????????????????????:
        _16376_ = b[247:240];
      64'b????????????????????????????????1???????????????????????????????:
        _16376_ = b[255:248];
      64'b???????????????????????????????1????????????????????????????????:
        _16376_ = b[263:256];
      64'b??????????????????????????????1?????????????????????????????????:
        _16376_ = b[271:264];
      64'b?????????????????????????????1??????????????????????????????????:
        _16376_ = b[279:272];
      64'b????????????????????????????1???????????????????????????????????:
        _16376_ = b[287:280];
      64'b???????????????????????????1????????????????????????????????????:
        _16376_ = b[295:288];
      64'b??????????????????????????1?????????????????????????????????????:
        _16376_ = b[303:296];
      64'b?????????????????????????1??????????????????????????????????????:
        _16376_ = b[311:304];
      64'b????????????????????????1???????????????????????????????????????:
        _16376_ = b[319:312];
      64'b???????????????????????1????????????????????????????????????????:
        _16376_ = b[327:320];
      64'b??????????????????????1?????????????????????????????????????????:
        _16376_ = b[335:328];
      64'b?????????????????????1??????????????????????????????????????????:
        _16376_ = b[343:336];
      64'b????????????????????1???????????????????????????????????????????:
        _16376_ = b[351:344];
      64'b???????????????????1????????????????????????????????????????????:
        _16376_ = b[359:352];
      64'b??????????????????1?????????????????????????????????????????????:
        _16376_ = b[367:360];
      64'b?????????????????1??????????????????????????????????????????????:
        _16376_ = b[375:368];
      64'b????????????????1???????????????????????????????????????????????:
        _16376_ = b[383:376];
      64'b???????????????1????????????????????????????????????????????????:
        _16376_ = b[391:384];
      64'b??????????????1?????????????????????????????????????????????????:
        _16376_ = b[399:392];
      64'b?????????????1??????????????????????????????????????????????????:
        _16376_ = b[407:400];
      64'b????????????1???????????????????????????????????????????????????:
        _16376_ = b[415:408];
      64'b???????????1????????????????????????????????????????????????????:
        _16376_ = b[423:416];
      64'b??????????1?????????????????????????????????????????????????????:
        _16376_ = b[431:424];
      64'b?????????1??????????????????????????????????????????????????????:
        _16376_ = b[439:432];
      64'b????????1???????????????????????????????????????????????????????:
        _16376_ = b[447:440];
      64'b???????1????????????????????????????????????????????????????????:
        _16376_ = b[455:448];
      64'b??????1?????????????????????????????????????????????????????????:
        _16376_ = b[463:456];
      64'b?????1??????????????????????????????????????????????????????????:
        _16376_ = b[471:464];
      64'b????1???????????????????????????????????????????????????????????:
        _16376_ = b[479:472];
      64'b???1????????????????????????????????????????????????????????????:
        _16376_ = b[487:480];
      64'b??1?????????????????????????????????????????????????????????????:
        _16376_ = b[495:488];
      64'b?1??????????????????????????????????????????????????????????????:
        _16376_ = b[503:496];
      64'b1???????????????????????????????????????????????????????????????:
        _16376_ = b[511:504];
      default:
        _16376_ = a;
    endcase
  endfunction
  assign vec_data_063 = _16376_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496], data_d1[511:504] }, { _06985_, _06984_, _06983_, _06982_, _06981_, _06980_, _06979_, _06978_, _06977_, _06976_, _06975_, _06974_, _06973_, _06972_, _06971_, _06970_, _06969_, _06968_, _06967_, _06966_, _06965_, _06964_, _06963_, _06962_, _06961_, _06960_, _06959_, _06958_, _06957_, _06956_, _06955_, _06954_, _06953_, _06952_, _06951_, _06950_, _06949_, _06948_, _06947_, _06946_, _06945_, _06944_, _06943_, _06942_, _06941_, _06940_, _06939_, _06938_, _06937_, _06936_, _06935_, _06934_, _06933_, _06932_, _06931_, _06930_, _06929_, _06928_, _06927_, _06926_, _06925_, _06924_, _06923_, _06922_ });
  assign _06922_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 7'b1000000;
  assign _06923_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111111;
  assign _06924_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111110;
  assign _06925_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111101;
  assign _06926_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111100;
  assign _06927_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111011;
  assign _06928_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111010;
  assign _06929_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111001;
  assign _06930_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b111000;
  assign _06931_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110111;
  assign _06932_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110110;
  assign _06933_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110101;
  assign _06934_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110100;
  assign _06935_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110011;
  assign _06936_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110010;
  assign _06937_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110001;
  assign _06938_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b110000;
  assign _06939_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101111;
  assign _06940_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101110;
  assign _06941_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101101;
  assign _06942_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101100;
  assign _06943_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101011;
  assign _06944_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101010;
  assign _06945_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101001;
  assign _06946_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b101000;
  assign _06947_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6450|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100111;
  assign _06948_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6449|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100110;
  assign _06949_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6448|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100101;
  assign _06950_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6447|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100100;
  assign _06951_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6446|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100011;
  assign _06952_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6445|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100010;
  assign _06953_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6444|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100001;
  assign _06954_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 6'b100000;
  assign _06955_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11111;
  assign _06956_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11110;
  assign _06957_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11101;
  assign _06958_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11100;
  assign _06959_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11011;
  assign _06960_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11010;
  assign _06961_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11001;
  assign _06962_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b11000;
  assign _06963_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10111;
  assign _06964_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10110;
  assign _06965_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10101;
  assign _06966_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10100;
  assign _06967_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10011;
  assign _06968_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10010;
  assign _06969_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10001;
  assign _06970_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 5'b10000;
  assign _06971_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1111;
  assign _06972_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1110;
  assign _06973_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1101;
  assign _06974_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1100;
  assign _06975_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1011;
  assign _06976_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1010;
  assign _06977_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1001;
  assign _06978_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 4'b1000;
  assign _06979_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 3'b111;
  assign _06980_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 3'b110;
  assign _06981_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 3'b101;
  assign _06982_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 3'b100;
  assign _06983_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 2'b11;
  assign _06984_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 2'b10;
  assign _06985_ = vec_sum_063_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6411" *) 1'b1;
  function [7:0] _16441_;
    input [7:0] a;
    input [503:0] b;
    input [62:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *)
    (* parallel_case *)
    casez (s)
      63'b??????????????????????????????????????????????????????????????1:
        _16441_ = b[7:0];
      63'b?????????????????????????????????????????????????????????????1?:
        _16441_ = b[15:8];
      63'b????????????????????????????????????????????????????????????1??:
        _16441_ = b[23:16];
      63'b???????????????????????????????????????????????????????????1???:
        _16441_ = b[31:24];
      63'b??????????????????????????????????????????????????????????1????:
        _16441_ = b[39:32];
      63'b?????????????????????????????????????????????????????????1?????:
        _16441_ = b[47:40];
      63'b????????????????????????????????????????????????????????1??????:
        _16441_ = b[55:48];
      63'b???????????????????????????????????????????????????????1???????:
        _16441_ = b[63:56];
      63'b??????????????????????????????????????????????????????1????????:
        _16441_ = b[71:64];
      63'b?????????????????????????????????????????????????????1?????????:
        _16441_ = b[79:72];
      63'b????????????????????????????????????????????????????1??????????:
        _16441_ = b[87:80];
      63'b???????????????????????????????????????????????????1???????????:
        _16441_ = b[95:88];
      63'b??????????????????????????????????????????????????1????????????:
        _16441_ = b[103:96];
      63'b?????????????????????????????????????????????????1?????????????:
        _16441_ = b[111:104];
      63'b????????????????????????????????????????????????1??????????????:
        _16441_ = b[119:112];
      63'b???????????????????????????????????????????????1???????????????:
        _16441_ = b[127:120];
      63'b??????????????????????????????????????????????1????????????????:
        _16441_ = b[135:128];
      63'b?????????????????????????????????????????????1?????????????????:
        _16441_ = b[143:136];
      63'b????????????????????????????????????????????1??????????????????:
        _16441_ = b[151:144];
      63'b???????????????????????????????????????????1???????????????????:
        _16441_ = b[159:152];
      63'b??????????????????????????????????????????1????????????????????:
        _16441_ = b[167:160];
      63'b?????????????????????????????????????????1?????????????????????:
        _16441_ = b[175:168];
      63'b????????????????????????????????????????1??????????????????????:
        _16441_ = b[183:176];
      63'b???????????????????????????????????????1???????????????????????:
        _16441_ = b[191:184];
      63'b??????????????????????????????????????1????????????????????????:
        _16441_ = b[199:192];
      63'b?????????????????????????????????????1?????????????????????????:
        _16441_ = b[207:200];
      63'b????????????????????????????????????1??????????????????????????:
        _16441_ = b[215:208];
      63'b???????????????????????????????????1???????????????????????????:
        _16441_ = b[223:216];
      63'b??????????????????????????????????1????????????????????????????:
        _16441_ = b[231:224];
      63'b?????????????????????????????????1?????????????????????????????:
        _16441_ = b[239:232];
      63'b????????????????????????????????1??????????????????????????????:
        _16441_ = b[247:240];
      63'b???????????????????????????????1???????????????????????????????:
        _16441_ = b[255:248];
      63'b??????????????????????????????1????????????????????????????????:
        _16441_ = b[263:256];
      63'b?????????????????????????????1?????????????????????????????????:
        _16441_ = b[271:264];
      63'b????????????????????????????1??????????????????????????????????:
        _16441_ = b[279:272];
      63'b???????????????????????????1???????????????????????????????????:
        _16441_ = b[287:280];
      63'b??????????????????????????1????????????????????????????????????:
        _16441_ = b[295:288];
      63'b?????????????????????????1?????????????????????????????????????:
        _16441_ = b[303:296];
      63'b????????????????????????1??????????????????????????????????????:
        _16441_ = b[311:304];
      63'b???????????????????????1???????????????????????????????????????:
        _16441_ = b[319:312];
      63'b??????????????????????1????????????????????????????????????????:
        _16441_ = b[327:320];
      63'b?????????????????????1?????????????????????????????????????????:
        _16441_ = b[335:328];
      63'b????????????????????1??????????????????????????????????????????:
        _16441_ = b[343:336];
      63'b???????????????????1???????????????????????????????????????????:
        _16441_ = b[351:344];
      63'b??????????????????1????????????????????????????????????????????:
        _16441_ = b[359:352];
      63'b?????????????????1?????????????????????????????????????????????:
        _16441_ = b[367:360];
      63'b????????????????1??????????????????????????????????????????????:
        _16441_ = b[375:368];
      63'b???????????????1???????????????????????????????????????????????:
        _16441_ = b[383:376];
      63'b??????????????1????????????????????????????????????????????????:
        _16441_ = b[391:384];
      63'b?????????????1?????????????????????????????????????????????????:
        _16441_ = b[399:392];
      63'b????????????1??????????????????????????????????????????????????:
        _16441_ = b[407:400];
      63'b???????????1???????????????????????????????????????????????????:
        _16441_ = b[415:408];
      63'b??????????1????????????????????????????????????????????????????:
        _16441_ = b[423:416];
      63'b?????????1?????????????????????????????????????????????????????:
        _16441_ = b[431:424];
      63'b????????1??????????????????????????????????????????????????????:
        _16441_ = b[439:432];
      63'b???????1???????????????????????????????????????????????????????:
        _16441_ = b[447:440];
      63'b??????1????????????????????????????????????????????????????????:
        _16441_ = b[455:448];
      63'b?????1?????????????????????????????????????????????????????????:
        _16441_ = b[463:456];
      63'b????1??????????????????????????????????????????????????????????:
        _16441_ = b[471:464];
      63'b???1???????????????????????????????????????????????????????????:
        _16441_ = b[479:472];
      63'b??1????????????????????????????????????????????????????????????:
        _16441_ = b[487:480];
      63'b?1?????????????????????????????????????????????????????????????:
        _16441_ = b[495:488];
      63'b1??????????????????????????????????????????????????????????????:
        _16441_ = b[503:496];
      default:
        _16441_ = a;
    endcase
  endfunction
  assign vec_data_062 = _16441_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488], data_d1[503:496] }, { _07048_, _07047_, _07046_, _07045_, _07044_, _07043_, _07042_, _07041_, _07040_, _07039_, _07038_, _07037_, _07036_, _07035_, _07034_, _07033_, _07032_, _07031_, _07030_, _07029_, _07028_, _07027_, _07026_, _07025_, _07024_, _07023_, _07022_, _07021_, _07020_, _07019_, _07018_, _07017_, _07016_, _07015_, _07014_, _07013_, _07012_, _07011_, _07010_, _07009_, _07008_, _07007_, _07006_, _07005_, _07004_, _07003_, _07002_, _07001_, _07000_, _06999_, _06998_, _06997_, _06996_, _06995_, _06994_, _06993_, _06992_, _06991_, _06990_, _06989_, _06988_, _06987_, _06986_ });
  assign _06986_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111111;
  assign _06987_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111110;
  assign _06988_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111101;
  assign _06989_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111100;
  assign _06990_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111011;
  assign _06991_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111010;
  assign _06992_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111001;
  assign _06993_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b111000;
  assign _06994_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110111;
  assign _06995_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110110;
  assign _06996_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110101;
  assign _06997_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110100;
  assign _06998_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110011;
  assign _06999_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110010;
  assign _07000_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110001;
  assign _07001_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b110000;
  assign _07002_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101111;
  assign _07003_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101110;
  assign _07004_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101101;
  assign _07005_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101100;
  assign _07006_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101011;
  assign _07007_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101010;
  assign _07008_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101001;
  assign _07009_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b101000;
  assign _07010_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100111;
  assign _07011_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100110;
  assign _07012_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100101;
  assign _07013_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100100;
  assign _07014_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100011;
  assign _07015_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100010;
  assign _07016_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100001;
  assign _07017_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 6'b100000;
  assign _07018_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11111;
  assign _07019_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11110;
  assign _07020_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11101;
  assign _07021_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11100;
  assign _07022_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11011;
  assign _07023_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11010;
  assign _07024_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11001;
  assign _07025_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b11000;
  assign _07026_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10111;
  assign _07027_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10110;
  assign _07028_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10101;
  assign _07029_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10100;
  assign _07030_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10011;
  assign _07031_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10010;
  assign _07032_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10001;
  assign _07033_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 5'b10000;
  assign _07034_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1111;
  assign _07035_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1110;
  assign _07036_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1101;
  assign _07037_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1100;
  assign _07038_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1011;
  assign _07039_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1010;
  assign _07040_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1001;
  assign _07041_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 4'b1000;
  assign _07042_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 3'b111;
  assign _07043_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 3'b110;
  assign _07044_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 3'b101;
  assign _07045_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 3'b100;
  assign _07046_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 2'b11;
  assign _07047_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 2'b10;
  assign _07048_ = vec_sum_062_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6340" *) 1'b1;
  function [7:0] _16505_;
    input [7:0] a;
    input [495:0] b;
    input [61:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *)
    (* parallel_case *)
    casez (s)
      62'b?????????????????????????????????????????????????????????????1:
        _16505_ = b[7:0];
      62'b????????????????????????????????????????????????????????????1?:
        _16505_ = b[15:8];
      62'b???????????????????????????????????????????????????????????1??:
        _16505_ = b[23:16];
      62'b??????????????????????????????????????????????????????????1???:
        _16505_ = b[31:24];
      62'b?????????????????????????????????????????????????????????1????:
        _16505_ = b[39:32];
      62'b????????????????????????????????????????????????????????1?????:
        _16505_ = b[47:40];
      62'b???????????????????????????????????????????????????????1??????:
        _16505_ = b[55:48];
      62'b??????????????????????????????????????????????????????1???????:
        _16505_ = b[63:56];
      62'b?????????????????????????????????????????????????????1????????:
        _16505_ = b[71:64];
      62'b????????????????????????????????????????????????????1?????????:
        _16505_ = b[79:72];
      62'b???????????????????????????????????????????????????1??????????:
        _16505_ = b[87:80];
      62'b??????????????????????????????????????????????????1???????????:
        _16505_ = b[95:88];
      62'b?????????????????????????????????????????????????1????????????:
        _16505_ = b[103:96];
      62'b????????????????????????????????????????????????1?????????????:
        _16505_ = b[111:104];
      62'b???????????????????????????????????????????????1??????????????:
        _16505_ = b[119:112];
      62'b??????????????????????????????????????????????1???????????????:
        _16505_ = b[127:120];
      62'b?????????????????????????????????????????????1????????????????:
        _16505_ = b[135:128];
      62'b????????????????????????????????????????????1?????????????????:
        _16505_ = b[143:136];
      62'b???????????????????????????????????????????1??????????????????:
        _16505_ = b[151:144];
      62'b??????????????????????????????????????????1???????????????????:
        _16505_ = b[159:152];
      62'b?????????????????????????????????????????1????????????????????:
        _16505_ = b[167:160];
      62'b????????????????????????????????????????1?????????????????????:
        _16505_ = b[175:168];
      62'b???????????????????????????????????????1??????????????????????:
        _16505_ = b[183:176];
      62'b??????????????????????????????????????1???????????????????????:
        _16505_ = b[191:184];
      62'b?????????????????????????????????????1????????????????????????:
        _16505_ = b[199:192];
      62'b????????????????????????????????????1?????????????????????????:
        _16505_ = b[207:200];
      62'b???????????????????????????????????1??????????????????????????:
        _16505_ = b[215:208];
      62'b??????????????????????????????????1???????????????????????????:
        _16505_ = b[223:216];
      62'b?????????????????????????????????1????????????????????????????:
        _16505_ = b[231:224];
      62'b????????????????????????????????1?????????????????????????????:
        _16505_ = b[239:232];
      62'b???????????????????????????????1??????????????????????????????:
        _16505_ = b[247:240];
      62'b??????????????????????????????1???????????????????????????????:
        _16505_ = b[255:248];
      62'b?????????????????????????????1????????????????????????????????:
        _16505_ = b[263:256];
      62'b????????????????????????????1?????????????????????????????????:
        _16505_ = b[271:264];
      62'b???????????????????????????1??????????????????????????????????:
        _16505_ = b[279:272];
      62'b??????????????????????????1???????????????????????????????????:
        _16505_ = b[287:280];
      62'b?????????????????????????1????????????????????????????????????:
        _16505_ = b[295:288];
      62'b????????????????????????1?????????????????????????????????????:
        _16505_ = b[303:296];
      62'b???????????????????????1??????????????????????????????????????:
        _16505_ = b[311:304];
      62'b??????????????????????1???????????????????????????????????????:
        _16505_ = b[319:312];
      62'b?????????????????????1????????????????????????????????????????:
        _16505_ = b[327:320];
      62'b????????????????????1?????????????????????????????????????????:
        _16505_ = b[335:328];
      62'b???????????????????1??????????????????????????????????????????:
        _16505_ = b[343:336];
      62'b??????????????????1???????????????????????????????????????????:
        _16505_ = b[351:344];
      62'b?????????????????1????????????????????????????????????????????:
        _16505_ = b[359:352];
      62'b????????????????1?????????????????????????????????????????????:
        _16505_ = b[367:360];
      62'b???????????????1??????????????????????????????????????????????:
        _16505_ = b[375:368];
      62'b??????????????1???????????????????????????????????????????????:
        _16505_ = b[383:376];
      62'b?????????????1????????????????????????????????????????????????:
        _16505_ = b[391:384];
      62'b????????????1?????????????????????????????????????????????????:
        _16505_ = b[399:392];
      62'b???????????1??????????????????????????????????????????????????:
        _16505_ = b[407:400];
      62'b??????????1???????????????????????????????????????????????????:
        _16505_ = b[415:408];
      62'b?????????1????????????????????????????????????????????????????:
        _16505_ = b[423:416];
      62'b????????1?????????????????????????????????????????????????????:
        _16505_ = b[431:424];
      62'b???????1??????????????????????????????????????????????????????:
        _16505_ = b[439:432];
      62'b??????1???????????????????????????????????????????????????????:
        _16505_ = b[447:440];
      62'b?????1????????????????????????????????????????????????????????:
        _16505_ = b[455:448];
      62'b????1?????????????????????????????????????????????????????????:
        _16505_ = b[463:456];
      62'b???1??????????????????????????????????????????????????????????:
        _16505_ = b[471:464];
      62'b??1???????????????????????????????????????????????????????????:
        _16505_ = b[479:472];
      62'b?1????????????????????????????????????????????????????????????:
        _16505_ = b[487:480];
      62'b1?????????????????????????????????????????????????????????????:
        _16505_ = b[495:488];
      default:
        _16505_ = a;
    endcase
  endfunction
  assign vec_data_061 = _16505_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480], data_d1[495:488] }, { _07110_, _07109_, _07108_, _07107_, _07106_, _07105_, _07104_, _07103_, _07102_, _07101_, _07100_, _07099_, _07098_, _07097_, _07096_, _07095_, _07094_, _07093_, _07092_, _07091_, _07090_, _07089_, _07088_, _07087_, _07086_, _07085_, _07084_, _07083_, _07082_, _07081_, _07080_, _07079_, _07078_, _07077_, _07076_, _07075_, _07074_, _07073_, _07072_, _07071_, _07070_, _07069_, _07068_, _07067_, _07066_, _07065_, _07064_, _07063_, _07062_, _07061_, _07060_, _07059_, _07058_, _07057_, _07056_, _07055_, _07054_, _07053_, _07052_, _07051_, _07050_, _07049_ });
  assign _07049_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111110;
  assign _07050_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111101;
  assign _07051_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111100;
  assign _07052_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111011;
  assign _07053_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111010;
  assign _07054_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111001;
  assign _07055_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b111000;
  assign _07056_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110111;
  assign _07057_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110110;
  assign _07058_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110101;
  assign _07059_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110100;
  assign _07060_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110011;
  assign _07061_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110010;
  assign _07062_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110001;
  assign _07063_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b110000;
  assign _07064_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101111;
  assign _07065_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101110;
  assign _07066_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101101;
  assign _07067_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101100;
  assign _07068_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101011;
  assign _07069_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101010;
  assign _07070_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101001;
  assign _07071_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b101000;
  assign _07072_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100111;
  assign _07073_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100110;
  assign _07074_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100101;
  assign _07075_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100100;
  assign _07076_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100011;
  assign _07077_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100010;
  assign _07078_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100001;
  assign _07079_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 6'b100000;
  assign _07080_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11111;
  assign _07081_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11110;
  assign _07082_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11101;
  assign _07083_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11100;
  assign _07084_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11011;
  assign _07085_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11010;
  assign _07086_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11001;
  assign _07087_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b11000;
  assign _07088_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10111;
  assign _07089_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10110;
  assign _07090_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10101;
  assign _07091_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10100;
  assign _07092_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10011;
  assign _07093_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10010;
  assign _07094_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10001;
  assign _07095_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6286|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 5'b10000;
  assign _07096_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6285|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1111;
  assign _07097_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6284|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1110;
  assign _07098_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6283|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1101;
  assign _07099_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1100;
  assign _07100_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1011;
  assign _07101_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1010;
  assign _07102_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1001;
  assign _07103_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 4'b1000;
  assign _07104_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 3'b111;
  assign _07105_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 3'b110;
  assign _07106_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 3'b101;
  assign _07107_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 3'b100;
  assign _07108_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 2'b11;
  assign _07109_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 2'b10;
  assign _07110_ = vec_sum_061_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6270" *) 1'b1;
  function [7:0] _16568_;
    input [7:0] a;
    input [487:0] b;
    input [60:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *)
    (* parallel_case *)
    casez (s)
      61'b????????????????????????????????????????????????????????????1:
        _16568_ = b[7:0];
      61'b???????????????????????????????????????????????????????????1?:
        _16568_ = b[15:8];
      61'b??????????????????????????????????????????????????????????1??:
        _16568_ = b[23:16];
      61'b?????????????????????????????????????????????????????????1???:
        _16568_ = b[31:24];
      61'b????????????????????????????????????????????????????????1????:
        _16568_ = b[39:32];
      61'b???????????????????????????????????????????????????????1?????:
        _16568_ = b[47:40];
      61'b??????????????????????????????????????????????????????1??????:
        _16568_ = b[55:48];
      61'b?????????????????????????????????????????????????????1???????:
        _16568_ = b[63:56];
      61'b????????????????????????????????????????????????????1????????:
        _16568_ = b[71:64];
      61'b???????????????????????????????????????????????????1?????????:
        _16568_ = b[79:72];
      61'b??????????????????????????????????????????????????1??????????:
        _16568_ = b[87:80];
      61'b?????????????????????????????????????????????????1???????????:
        _16568_ = b[95:88];
      61'b????????????????????????????????????????????????1????????????:
        _16568_ = b[103:96];
      61'b???????????????????????????????????????????????1?????????????:
        _16568_ = b[111:104];
      61'b??????????????????????????????????????????????1??????????????:
        _16568_ = b[119:112];
      61'b?????????????????????????????????????????????1???????????????:
        _16568_ = b[127:120];
      61'b????????????????????????????????????????????1????????????????:
        _16568_ = b[135:128];
      61'b???????????????????????????????????????????1?????????????????:
        _16568_ = b[143:136];
      61'b??????????????????????????????????????????1??????????????????:
        _16568_ = b[151:144];
      61'b?????????????????????????????????????????1???????????????????:
        _16568_ = b[159:152];
      61'b????????????????????????????????????????1????????????????????:
        _16568_ = b[167:160];
      61'b???????????????????????????????????????1?????????????????????:
        _16568_ = b[175:168];
      61'b??????????????????????????????????????1??????????????????????:
        _16568_ = b[183:176];
      61'b?????????????????????????????????????1???????????????????????:
        _16568_ = b[191:184];
      61'b????????????????????????????????????1????????????????????????:
        _16568_ = b[199:192];
      61'b???????????????????????????????????1?????????????????????????:
        _16568_ = b[207:200];
      61'b??????????????????????????????????1??????????????????????????:
        _16568_ = b[215:208];
      61'b?????????????????????????????????1???????????????????????????:
        _16568_ = b[223:216];
      61'b????????????????????????????????1????????????????????????????:
        _16568_ = b[231:224];
      61'b???????????????????????????????1?????????????????????????????:
        _16568_ = b[239:232];
      61'b??????????????????????????????1??????????????????????????????:
        _16568_ = b[247:240];
      61'b?????????????????????????????1???????????????????????????????:
        _16568_ = b[255:248];
      61'b????????????????????????????1????????????????????????????????:
        _16568_ = b[263:256];
      61'b???????????????????????????1?????????????????????????????????:
        _16568_ = b[271:264];
      61'b??????????????????????????1??????????????????????????????????:
        _16568_ = b[279:272];
      61'b?????????????????????????1???????????????????????????????????:
        _16568_ = b[287:280];
      61'b????????????????????????1????????????????????????????????????:
        _16568_ = b[295:288];
      61'b???????????????????????1?????????????????????????????????????:
        _16568_ = b[303:296];
      61'b??????????????????????1??????????????????????????????????????:
        _16568_ = b[311:304];
      61'b?????????????????????1???????????????????????????????????????:
        _16568_ = b[319:312];
      61'b????????????????????1????????????????????????????????????????:
        _16568_ = b[327:320];
      61'b???????????????????1?????????????????????????????????????????:
        _16568_ = b[335:328];
      61'b??????????????????1??????????????????????????????????????????:
        _16568_ = b[343:336];
      61'b?????????????????1???????????????????????????????????????????:
        _16568_ = b[351:344];
      61'b????????????????1????????????????????????????????????????????:
        _16568_ = b[359:352];
      61'b???????????????1?????????????????????????????????????????????:
        _16568_ = b[367:360];
      61'b??????????????1??????????????????????????????????????????????:
        _16568_ = b[375:368];
      61'b?????????????1???????????????????????????????????????????????:
        _16568_ = b[383:376];
      61'b????????????1????????????????????????????????????????????????:
        _16568_ = b[391:384];
      61'b???????????1?????????????????????????????????????????????????:
        _16568_ = b[399:392];
      61'b??????????1??????????????????????????????????????????????????:
        _16568_ = b[407:400];
      61'b?????????1???????????????????????????????????????????????????:
        _16568_ = b[415:408];
      61'b????????1????????????????????????????????????????????????????:
        _16568_ = b[423:416];
      61'b???????1?????????????????????????????????????????????????????:
        _16568_ = b[431:424];
      61'b??????1??????????????????????????????????????????????????????:
        _16568_ = b[439:432];
      61'b?????1???????????????????????????????????????????????????????:
        _16568_ = b[447:440];
      61'b????1????????????????????????????????????????????????????????:
        _16568_ = b[455:448];
      61'b???1?????????????????????????????????????????????????????????:
        _16568_ = b[463:456];
      61'b??1??????????????????????????????????????????????????????????:
        _16568_ = b[471:464];
      61'b?1???????????????????????????????????????????????????????????:
        _16568_ = b[479:472];
      61'b1????????????????????????????????????????????????????????????:
        _16568_ = b[487:480];
      default:
        _16568_ = a;
    endcase
  endfunction
  assign vec_data_060 = _16568_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472], data_d1[487:480] }, { _07171_, _07170_, _07169_, _07168_, _07167_, _07166_, _07165_, _07164_, _07163_, _07162_, _07161_, _07160_, _07159_, _07158_, _07157_, _07156_, _07155_, _07154_, _07153_, _07152_, _07151_, _07150_, _07149_, _07148_, _07147_, _07146_, _07145_, _07144_, _07143_, _07142_, _07141_, _07140_, _07139_, _07138_, _07137_, _07136_, _07135_, _07134_, _07133_, _07132_, _07131_, _07130_, _07129_, _07128_, _07127_, _07126_, _07125_, _07124_, _07123_, _07122_, _07121_, _07120_, _07119_, _07118_, _07117_, _07116_, _07115_, _07114_, _07113_, _07112_, _07111_ });
  assign _07111_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111101;
  assign _07112_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111100;
  assign _07113_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111011;
  assign _07114_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111010;
  assign _07115_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111001;
  assign _07116_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b111000;
  assign _07117_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110111;
  assign _07118_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110110;
  assign _07119_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110101;
  assign _07120_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110100;
  assign _07121_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110011;
  assign _07122_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110010;
  assign _07123_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110001;
  assign _07124_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b110000;
  assign _07125_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101111;
  assign _07126_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101110;
  assign _07127_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101101;
  assign _07128_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101100;
  assign _07129_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101011;
  assign _07130_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101010;
  assign _07131_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101001;
  assign _07132_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b101000;
  assign _07133_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100111;
  assign _07134_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100110;
  assign _07135_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100101;
  assign _07136_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100100;
  assign _07137_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100011;
  assign _07138_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100010;
  assign _07139_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100001;
  assign _07140_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6233|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 6'b100000;
  assign _07141_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6232|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11111;
  assign _07142_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6231|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11110;
  assign _07143_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6230|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11101;
  assign _07144_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6229|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11100;
  assign _07145_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6228|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11011;
  assign _07146_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6227|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11010;
  assign _07147_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6226|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11001;
  assign _07148_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b11000;
  assign _07149_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10111;
  assign _07150_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10110;
  assign _07151_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10101;
  assign _07152_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10100;
  assign _07153_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10011;
  assign _07154_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10010;
  assign _07155_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10001;
  assign _07156_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 5'b10000;
  assign _07157_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1111;
  assign _07158_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1110;
  assign _07159_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1101;
  assign _07160_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1100;
  assign _07161_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1011;
  assign _07162_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1010;
  assign _07163_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1001;
  assign _07164_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 4'b1000;
  assign _07165_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 3'b111;
  assign _07166_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 3'b110;
  assign _07167_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 3'b101;
  assign _07168_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 3'b100;
  assign _07169_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 2'b11;
  assign _07170_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 2'b10;
  assign _07171_ = vec_sum_060_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6201" *) 1'b1;
  function [7:0] _16630_;
    input [7:0] a;
    input [479:0] b;
    input [59:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *)
    (* parallel_case *)
    casez (s)
      60'b???????????????????????????????????????????????????????????1:
        _16630_ = b[7:0];
      60'b??????????????????????????????????????????????????????????1?:
        _16630_ = b[15:8];
      60'b?????????????????????????????????????????????????????????1??:
        _16630_ = b[23:16];
      60'b????????????????????????????????????????????????????????1???:
        _16630_ = b[31:24];
      60'b???????????????????????????????????????????????????????1????:
        _16630_ = b[39:32];
      60'b??????????????????????????????????????????????????????1?????:
        _16630_ = b[47:40];
      60'b?????????????????????????????????????????????????????1??????:
        _16630_ = b[55:48];
      60'b????????????????????????????????????????????????????1???????:
        _16630_ = b[63:56];
      60'b???????????????????????????????????????????????????1????????:
        _16630_ = b[71:64];
      60'b??????????????????????????????????????????????????1?????????:
        _16630_ = b[79:72];
      60'b?????????????????????????????????????????????????1??????????:
        _16630_ = b[87:80];
      60'b????????????????????????????????????????????????1???????????:
        _16630_ = b[95:88];
      60'b???????????????????????????????????????????????1????????????:
        _16630_ = b[103:96];
      60'b??????????????????????????????????????????????1?????????????:
        _16630_ = b[111:104];
      60'b?????????????????????????????????????????????1??????????????:
        _16630_ = b[119:112];
      60'b????????????????????????????????????????????1???????????????:
        _16630_ = b[127:120];
      60'b???????????????????????????????????????????1????????????????:
        _16630_ = b[135:128];
      60'b??????????????????????????????????????????1?????????????????:
        _16630_ = b[143:136];
      60'b?????????????????????????????????????????1??????????????????:
        _16630_ = b[151:144];
      60'b????????????????????????????????????????1???????????????????:
        _16630_ = b[159:152];
      60'b???????????????????????????????????????1????????????????????:
        _16630_ = b[167:160];
      60'b??????????????????????????????????????1?????????????????????:
        _16630_ = b[175:168];
      60'b?????????????????????????????????????1??????????????????????:
        _16630_ = b[183:176];
      60'b????????????????????????????????????1???????????????????????:
        _16630_ = b[191:184];
      60'b???????????????????????????????????1????????????????????????:
        _16630_ = b[199:192];
      60'b??????????????????????????????????1?????????????????????????:
        _16630_ = b[207:200];
      60'b?????????????????????????????????1??????????????????????????:
        _16630_ = b[215:208];
      60'b????????????????????????????????1???????????????????????????:
        _16630_ = b[223:216];
      60'b???????????????????????????????1????????????????????????????:
        _16630_ = b[231:224];
      60'b??????????????????????????????1?????????????????????????????:
        _16630_ = b[239:232];
      60'b?????????????????????????????1??????????????????????????????:
        _16630_ = b[247:240];
      60'b????????????????????????????1???????????????????????????????:
        _16630_ = b[255:248];
      60'b???????????????????????????1????????????????????????????????:
        _16630_ = b[263:256];
      60'b??????????????????????????1?????????????????????????????????:
        _16630_ = b[271:264];
      60'b?????????????????????????1??????????????????????????????????:
        _16630_ = b[279:272];
      60'b????????????????????????1???????????????????????????????????:
        _16630_ = b[287:280];
      60'b???????????????????????1????????????????????????????????????:
        _16630_ = b[295:288];
      60'b??????????????????????1?????????????????????????????????????:
        _16630_ = b[303:296];
      60'b?????????????????????1??????????????????????????????????????:
        _16630_ = b[311:304];
      60'b????????????????????1???????????????????????????????????????:
        _16630_ = b[319:312];
      60'b???????????????????1????????????????????????????????????????:
        _16630_ = b[327:320];
      60'b??????????????????1?????????????????????????????????????????:
        _16630_ = b[335:328];
      60'b?????????????????1??????????????????????????????????????????:
        _16630_ = b[343:336];
      60'b????????????????1???????????????????????????????????????????:
        _16630_ = b[351:344];
      60'b???????????????1????????????????????????????????????????????:
        _16630_ = b[359:352];
      60'b??????????????1?????????????????????????????????????????????:
        _16630_ = b[367:360];
      60'b?????????????1??????????????????????????????????????????????:
        _16630_ = b[375:368];
      60'b????????????1???????????????????????????????????????????????:
        _16630_ = b[383:376];
      60'b???????????1????????????????????????????????????????????????:
        _16630_ = b[391:384];
      60'b??????????1?????????????????????????????????????????????????:
        _16630_ = b[399:392];
      60'b?????????1??????????????????????????????????????????????????:
        _16630_ = b[407:400];
      60'b????????1???????????????????????????????????????????????????:
        _16630_ = b[415:408];
      60'b???????1????????????????????????????????????????????????????:
        _16630_ = b[423:416];
      60'b??????1?????????????????????????????????????????????????????:
        _16630_ = b[431:424];
      60'b?????1??????????????????????????????????????????????????????:
        _16630_ = b[439:432];
      60'b????1???????????????????????????????????????????????????????:
        _16630_ = b[447:440];
      60'b???1????????????????????????????????????????????????????????:
        _16630_ = b[455:448];
      60'b??1?????????????????????????????????????????????????????????:
        _16630_ = b[463:456];
      60'b?1??????????????????????????????????????????????????????????:
        _16630_ = b[471:464];
      60'b1???????????????????????????????????????????????????????????:
        _16630_ = b[479:472];
      default:
        _16630_ = a;
    endcase
  endfunction
  assign vec_data_059 = _16630_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464], data_d1[479:472] }, { _07231_, _07230_, _07229_, _07228_, _07227_, _07226_, _07225_, _07224_, _07223_, _07222_, _07221_, _07220_, _07219_, _07218_, _07217_, _07216_, _07215_, _07214_, _07213_, _07212_, _07211_, _07210_, _07209_, _07208_, _07207_, _07206_, _07205_, _07204_, _07203_, _07202_, _07201_, _07200_, _07199_, _07198_, _07197_, _07196_, _07195_, _07194_, _07193_, _07192_, _07191_, _07190_, _07189_, _07188_, _07187_, _07186_, _07185_, _07184_, _07183_, _07182_, _07181_, _07180_, _07179_, _07178_, _07177_, _07176_, _07175_, _07174_, _07173_, _07172_ });
  assign _07172_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b111100;
  assign _07173_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b111011;
  assign _07174_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b111010;
  assign _07175_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b111001;
  assign _07176_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b111000;
  assign _07177_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110111;
  assign _07178_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110110;
  assign _07179_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110101;
  assign _07180_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110100;
  assign _07181_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110011;
  assign _07182_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110010;
  assign _07183_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110001;
  assign _07184_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b110000;
  assign _07185_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6180|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101111;
  assign _07186_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6179|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101110;
  assign _07187_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6178|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101101;
  assign _07188_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6177|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101100;
  assign _07189_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6176|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101011;
  assign _07190_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6175|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101010;
  assign _07191_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6174|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101001;
  assign _07192_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b101000;
  assign _07193_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100111;
  assign _07194_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100110;
  assign _07195_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100101;
  assign _07196_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100100;
  assign _07197_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100011;
  assign _07198_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100010;
  assign _07199_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100001;
  assign _07200_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 6'b100000;
  assign _07201_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11111;
  assign _07202_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11110;
  assign _07203_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11101;
  assign _07204_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11100;
  assign _07205_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11011;
  assign _07206_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11010;
  assign _07207_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11001;
  assign _07208_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b11000;
  assign _07209_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10111;
  assign _07210_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10110;
  assign _07211_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10101;
  assign _07212_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10100;
  assign _07213_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10011;
  assign _07214_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10010;
  assign _07215_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10001;
  assign _07216_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 5'b10000;
  assign _07217_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1111;
  assign _07218_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1110;
  assign _07219_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1101;
  assign _07220_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1100;
  assign _07221_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1011;
  assign _07222_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1010;
  assign _07223_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1001;
  assign _07224_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 4'b1000;
  assign _07225_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 3'b111;
  assign _07226_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 3'b110;
  assign _07227_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 3'b101;
  assign _07228_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 3'b100;
  assign _07229_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 2'b11;
  assign _07230_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 2'b10;
  assign _07231_ = vec_sum_059_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6133" *) 1'b1;
  function [7:0] _16691_;
    input [7:0] a;
    input [471:0] b;
    input [58:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *)
    (* parallel_case *)
    casez (s)
      59'b??????????????????????????????????????????????????????????1:
        _16691_ = b[7:0];
      59'b?????????????????????????????????????????????????????????1?:
        _16691_ = b[15:8];
      59'b????????????????????????????????????????????????????????1??:
        _16691_ = b[23:16];
      59'b???????????????????????????????????????????????????????1???:
        _16691_ = b[31:24];
      59'b??????????????????????????????????????????????????????1????:
        _16691_ = b[39:32];
      59'b?????????????????????????????????????????????????????1?????:
        _16691_ = b[47:40];
      59'b????????????????????????????????????????????????????1??????:
        _16691_ = b[55:48];
      59'b???????????????????????????????????????????????????1???????:
        _16691_ = b[63:56];
      59'b??????????????????????????????????????????????????1????????:
        _16691_ = b[71:64];
      59'b?????????????????????????????????????????????????1?????????:
        _16691_ = b[79:72];
      59'b????????????????????????????????????????????????1??????????:
        _16691_ = b[87:80];
      59'b???????????????????????????????????????????????1???????????:
        _16691_ = b[95:88];
      59'b??????????????????????????????????????????????1????????????:
        _16691_ = b[103:96];
      59'b?????????????????????????????????????????????1?????????????:
        _16691_ = b[111:104];
      59'b????????????????????????????????????????????1??????????????:
        _16691_ = b[119:112];
      59'b???????????????????????????????????????????1???????????????:
        _16691_ = b[127:120];
      59'b??????????????????????????????????????????1????????????????:
        _16691_ = b[135:128];
      59'b?????????????????????????????????????????1?????????????????:
        _16691_ = b[143:136];
      59'b????????????????????????????????????????1??????????????????:
        _16691_ = b[151:144];
      59'b???????????????????????????????????????1???????????????????:
        _16691_ = b[159:152];
      59'b??????????????????????????????????????1????????????????????:
        _16691_ = b[167:160];
      59'b?????????????????????????????????????1?????????????????????:
        _16691_ = b[175:168];
      59'b????????????????????????????????????1??????????????????????:
        _16691_ = b[183:176];
      59'b???????????????????????????????????1???????????????????????:
        _16691_ = b[191:184];
      59'b??????????????????????????????????1????????????????????????:
        _16691_ = b[199:192];
      59'b?????????????????????????????????1?????????????????????????:
        _16691_ = b[207:200];
      59'b????????????????????????????????1??????????????????????????:
        _16691_ = b[215:208];
      59'b???????????????????????????????1???????????????????????????:
        _16691_ = b[223:216];
      59'b??????????????????????????????1????????????????????????????:
        _16691_ = b[231:224];
      59'b?????????????????????????????1?????????????????????????????:
        _16691_ = b[239:232];
      59'b????????????????????????????1??????????????????????????????:
        _16691_ = b[247:240];
      59'b???????????????????????????1???????????????????????????????:
        _16691_ = b[255:248];
      59'b??????????????????????????1????????????????????????????????:
        _16691_ = b[263:256];
      59'b?????????????????????????1?????????????????????????????????:
        _16691_ = b[271:264];
      59'b????????????????????????1??????????????????????????????????:
        _16691_ = b[279:272];
      59'b???????????????????????1???????????????????????????????????:
        _16691_ = b[287:280];
      59'b??????????????????????1????????????????????????????????????:
        _16691_ = b[295:288];
      59'b?????????????????????1?????????????????????????????????????:
        _16691_ = b[303:296];
      59'b????????????????????1??????????????????????????????????????:
        _16691_ = b[311:304];
      59'b???????????????????1???????????????????????????????????????:
        _16691_ = b[319:312];
      59'b??????????????????1????????????????????????????????????????:
        _16691_ = b[327:320];
      59'b?????????????????1?????????????????????????????????????????:
        _16691_ = b[335:328];
      59'b????????????????1??????????????????????????????????????????:
        _16691_ = b[343:336];
      59'b???????????????1???????????????????????????????????????????:
        _16691_ = b[351:344];
      59'b??????????????1????????????????????????????????????????????:
        _16691_ = b[359:352];
      59'b?????????????1?????????????????????????????????????????????:
        _16691_ = b[367:360];
      59'b????????????1??????????????????????????????????????????????:
        _16691_ = b[375:368];
      59'b???????????1???????????????????????????????????????????????:
        _16691_ = b[383:376];
      59'b??????????1????????????????????????????????????????????????:
        _16691_ = b[391:384];
      59'b?????????1?????????????????????????????????????????????????:
        _16691_ = b[399:392];
      59'b????????1??????????????????????????????????????????????????:
        _16691_ = b[407:400];
      59'b???????1???????????????????????????????????????????????????:
        _16691_ = b[415:408];
      59'b??????1????????????????????????????????????????????????????:
        _16691_ = b[423:416];
      59'b?????1?????????????????????????????????????????????????????:
        _16691_ = b[431:424];
      59'b????1??????????????????????????????????????????????????????:
        _16691_ = b[439:432];
      59'b???1???????????????????????????????????????????????????????:
        _16691_ = b[447:440];
      59'b??1????????????????????????????????????????????????????????:
        _16691_ = b[455:448];
      59'b?1?????????????????????????????????????????????????????????:
        _16691_ = b[463:456];
      59'b1??????????????????????????????????????????????????????????:
        _16691_ = b[471:464];
      default:
        _16691_ = a;
    endcase
  endfunction
  assign vec_data_058 = _16691_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456], data_d1[471:464] }, { _07290_, _07289_, _07288_, _07287_, _07286_, _07285_, _07284_, _07283_, _07282_, _07281_, _07280_, _07279_, _07278_, _07277_, _07276_, _07275_, _07274_, _07273_, _07272_, _07271_, _07270_, _07269_, _07268_, _07267_, _07266_, _07265_, _07264_, _07263_, _07262_, _07261_, _07260_, _07259_, _07258_, _07257_, _07256_, _07255_, _07254_, _07253_, _07252_, _07251_, _07250_, _07249_, _07248_, _07247_, _07246_, _07245_, _07244_, _07243_, _07242_, _07241_, _07240_, _07239_, _07238_, _07237_, _07236_, _07235_, _07234_, _07233_, _07232_ });
  assign _07232_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6125|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b111011;
  assign _07233_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6124|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b111010;
  assign _07234_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b111001;
  assign _07235_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b111000;
  assign _07236_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110111;
  assign _07237_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110110;
  assign _07238_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110101;
  assign _07239_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110100;
  assign _07240_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110011;
  assign _07241_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110010;
  assign _07242_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110001;
  assign _07243_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b110000;
  assign _07244_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101111;
  assign _07245_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101110;
  assign _07246_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101101;
  assign _07247_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101100;
  assign _07248_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101011;
  assign _07249_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101010;
  assign _07250_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101001;
  assign _07251_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b101000;
  assign _07252_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100111;
  assign _07253_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100110;
  assign _07254_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100101;
  assign _07255_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100100;
  assign _07256_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100011;
  assign _07257_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100010;
  assign _07258_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100001;
  assign _07259_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 6'b100000;
  assign _07260_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11111;
  assign _07261_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11110;
  assign _07262_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11101;
  assign _07263_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11100;
  assign _07264_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11011;
  assign _07265_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11010;
  assign _07266_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11001;
  assign _07267_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b11000;
  assign _07268_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10111;
  assign _07269_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10110;
  assign _07270_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10101;
  assign _07271_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10100;
  assign _07272_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10011;
  assign _07273_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10010;
  assign _07274_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10001;
  assign _07275_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 5'b10000;
  assign _07276_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1111;
  assign _07277_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6080|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1110;
  assign _07278_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6079|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1101;
  assign _07279_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1100;
  assign _07280_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1011;
  assign _07281_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1010;
  assign _07282_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1001;
  assign _07283_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 4'b1000;
  assign _07284_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 3'b111;
  assign _07285_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 3'b110;
  assign _07286_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 3'b101;
  assign _07287_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 3'b100;
  assign _07288_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 2'b11;
  assign _07289_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 2'b10;
  assign _07290_ = vec_sum_058_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6066" *) 1'b1;
  function [7:0] _16751_;
    input [7:0] a;
    input [463:0] b;
    input [57:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *)
    (* parallel_case *)
    casez (s)
      58'b?????????????????????????????????????????????????????????1:
        _16751_ = b[7:0];
      58'b????????????????????????????????????????????????????????1?:
        _16751_ = b[15:8];
      58'b???????????????????????????????????????????????????????1??:
        _16751_ = b[23:16];
      58'b??????????????????????????????????????????????????????1???:
        _16751_ = b[31:24];
      58'b?????????????????????????????????????????????????????1????:
        _16751_ = b[39:32];
      58'b????????????????????????????????????????????????????1?????:
        _16751_ = b[47:40];
      58'b???????????????????????????????????????????????????1??????:
        _16751_ = b[55:48];
      58'b??????????????????????????????????????????????????1???????:
        _16751_ = b[63:56];
      58'b?????????????????????????????????????????????????1????????:
        _16751_ = b[71:64];
      58'b????????????????????????????????????????????????1?????????:
        _16751_ = b[79:72];
      58'b???????????????????????????????????????????????1??????????:
        _16751_ = b[87:80];
      58'b??????????????????????????????????????????????1???????????:
        _16751_ = b[95:88];
      58'b?????????????????????????????????????????????1????????????:
        _16751_ = b[103:96];
      58'b????????????????????????????????????????????1?????????????:
        _16751_ = b[111:104];
      58'b???????????????????????????????????????????1??????????????:
        _16751_ = b[119:112];
      58'b??????????????????????????????????????????1???????????????:
        _16751_ = b[127:120];
      58'b?????????????????????????????????????????1????????????????:
        _16751_ = b[135:128];
      58'b????????????????????????????????????????1?????????????????:
        _16751_ = b[143:136];
      58'b???????????????????????????????????????1??????????????????:
        _16751_ = b[151:144];
      58'b??????????????????????????????????????1???????????????????:
        _16751_ = b[159:152];
      58'b?????????????????????????????????????1????????????????????:
        _16751_ = b[167:160];
      58'b????????????????????????????????????1?????????????????????:
        _16751_ = b[175:168];
      58'b???????????????????????????????????1??????????????????????:
        _16751_ = b[183:176];
      58'b??????????????????????????????????1???????????????????????:
        _16751_ = b[191:184];
      58'b?????????????????????????????????1????????????????????????:
        _16751_ = b[199:192];
      58'b????????????????????????????????1?????????????????????????:
        _16751_ = b[207:200];
      58'b???????????????????????????????1??????????????????????????:
        _16751_ = b[215:208];
      58'b??????????????????????????????1???????????????????????????:
        _16751_ = b[223:216];
      58'b?????????????????????????????1????????????????????????????:
        _16751_ = b[231:224];
      58'b????????????????????????????1?????????????????????????????:
        _16751_ = b[239:232];
      58'b???????????????????????????1??????????????????????????????:
        _16751_ = b[247:240];
      58'b??????????????????????????1???????????????????????????????:
        _16751_ = b[255:248];
      58'b?????????????????????????1????????????????????????????????:
        _16751_ = b[263:256];
      58'b????????????????????????1?????????????????????????????????:
        _16751_ = b[271:264];
      58'b???????????????????????1??????????????????????????????????:
        _16751_ = b[279:272];
      58'b??????????????????????1???????????????????????????????????:
        _16751_ = b[287:280];
      58'b?????????????????????1????????????????????????????????????:
        _16751_ = b[295:288];
      58'b????????????????????1?????????????????????????????????????:
        _16751_ = b[303:296];
      58'b???????????????????1??????????????????????????????????????:
        _16751_ = b[311:304];
      58'b??????????????????1???????????????????????????????????????:
        _16751_ = b[319:312];
      58'b?????????????????1????????????????????????????????????????:
        _16751_ = b[327:320];
      58'b????????????????1?????????????????????????????????????????:
        _16751_ = b[335:328];
      58'b???????????????1??????????????????????????????????????????:
        _16751_ = b[343:336];
      58'b??????????????1???????????????????????????????????????????:
        _16751_ = b[351:344];
      58'b?????????????1????????????????????????????????????????????:
        _16751_ = b[359:352];
      58'b????????????1?????????????????????????????????????????????:
        _16751_ = b[367:360];
      58'b???????????1??????????????????????????????????????????????:
        _16751_ = b[375:368];
      58'b??????????1???????????????????????????????????????????????:
        _16751_ = b[383:376];
      58'b?????????1????????????????????????????????????????????????:
        _16751_ = b[391:384];
      58'b????????1?????????????????????????????????????????????????:
        _16751_ = b[399:392];
      58'b???????1??????????????????????????????????????????????????:
        _16751_ = b[407:400];
      58'b??????1???????????????????????????????????????????????????:
        _16751_ = b[415:408];
      58'b?????1????????????????????????????????????????????????????:
        _16751_ = b[423:416];
      58'b????1?????????????????????????????????????????????????????:
        _16751_ = b[431:424];
      58'b???1??????????????????????????????????????????????????????:
        _16751_ = b[439:432];
      58'b??1???????????????????????????????????????????????????????:
        _16751_ = b[447:440];
      58'b?1????????????????????????????????????????????????????????:
        _16751_ = b[455:448];
      58'b1?????????????????????????????????????????????????????????:
        _16751_ = b[463:456];
      default:
        _16751_ = a;
    endcase
  endfunction
  assign vec_data_057 = _16751_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448], data_d1[463:456] }, { _07348_, _07347_, _07346_, _07345_, _07344_, _07343_, _07342_, _07341_, _07340_, _07339_, _07338_, _07337_, _07336_, _07335_, _07334_, _07333_, _07332_, _07331_, _07330_, _07329_, _07328_, _07327_, _07326_, _07325_, _07324_, _07323_, _07322_, _07321_, _07320_, _07319_, _07318_, _07317_, _07316_, _07315_, _07314_, _07313_, _07312_, _07311_, _07310_, _07309_, _07308_, _07307_, _07306_, _07305_, _07304_, _07303_, _07302_, _07301_, _07300_, _07299_, _07298_, _07297_, _07296_, _07295_, _07294_, _07293_, _07292_, _07291_ });
  assign _07291_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b111010;
  assign _07292_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b111001;
  assign _07293_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b111000;
  assign _07294_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110111;
  assign _07295_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110110;
  assign _07296_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110101;
  assign _07297_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110100;
  assign _07298_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110011;
  assign _07299_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110010;
  assign _07300_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110001;
  assign _07301_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b110000;
  assign _07302_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101111;
  assign _07303_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101110;
  assign _07304_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101101;
  assign _07305_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101100;
  assign _07306_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101011;
  assign _07307_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101010;
  assign _07308_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101001;
  assign _07309_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b101000;
  assign _07310_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100111;
  assign _07311_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100110;
  assign _07312_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100101;
  assign _07313_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100100;
  assign _07314_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100011;
  assign _07315_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100010;
  assign _07316_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100001;
  assign _07317_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 6'b100000;
  assign _07318_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11111;
  assign _07319_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11110;
  assign _07320_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11101;
  assign _07321_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11100;
  assign _07322_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11011;
  assign _07323_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6026|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11010;
  assign _07324_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6025|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11001;
  assign _07325_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6024|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b11000;
  assign _07326_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10111;
  assign _07327_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10110;
  assign _07328_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10101;
  assign _07329_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10100;
  assign _07330_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10011;
  assign _07331_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10010;
  assign _07332_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10001;
  assign _07333_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 5'b10000;
  assign _07334_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1111;
  assign _07335_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1110;
  assign _07336_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1101;
  assign _07337_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1100;
  assign _07338_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1011;
  assign _07339_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1010;
  assign _07340_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1001;
  assign _07341_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 4'b1000;
  assign _07342_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 3'b111;
  assign _07343_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 3'b110;
  assign _07344_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 3'b101;
  assign _07345_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 3'b100;
  assign _07346_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 2'b11;
  assign _07347_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 2'b10;
  assign _07348_ = vec_sum_057_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:6000" *) 1'b1;
  function [7:0] _16810_;
    input [7:0] a;
    input [455:0] b;
    input [56:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *)
    (* parallel_case *)
    casez (s)
      57'b????????????????????????????????????????????????????????1:
        _16810_ = b[7:0];
      57'b???????????????????????????????????????????????????????1?:
        _16810_ = b[15:8];
      57'b??????????????????????????????????????????????????????1??:
        _16810_ = b[23:16];
      57'b?????????????????????????????????????????????????????1???:
        _16810_ = b[31:24];
      57'b????????????????????????????????????????????????????1????:
        _16810_ = b[39:32];
      57'b???????????????????????????????????????????????????1?????:
        _16810_ = b[47:40];
      57'b??????????????????????????????????????????????????1??????:
        _16810_ = b[55:48];
      57'b?????????????????????????????????????????????????1???????:
        _16810_ = b[63:56];
      57'b????????????????????????????????????????????????1????????:
        _16810_ = b[71:64];
      57'b???????????????????????????????????????????????1?????????:
        _16810_ = b[79:72];
      57'b??????????????????????????????????????????????1??????????:
        _16810_ = b[87:80];
      57'b?????????????????????????????????????????????1???????????:
        _16810_ = b[95:88];
      57'b????????????????????????????????????????????1????????????:
        _16810_ = b[103:96];
      57'b???????????????????????????????????????????1?????????????:
        _16810_ = b[111:104];
      57'b??????????????????????????????????????????1??????????????:
        _16810_ = b[119:112];
      57'b?????????????????????????????????????????1???????????????:
        _16810_ = b[127:120];
      57'b????????????????????????????????????????1????????????????:
        _16810_ = b[135:128];
      57'b???????????????????????????????????????1?????????????????:
        _16810_ = b[143:136];
      57'b??????????????????????????????????????1??????????????????:
        _16810_ = b[151:144];
      57'b?????????????????????????????????????1???????????????????:
        _16810_ = b[159:152];
      57'b????????????????????????????????????1????????????????????:
        _16810_ = b[167:160];
      57'b???????????????????????????????????1?????????????????????:
        _16810_ = b[175:168];
      57'b??????????????????????????????????1??????????????????????:
        _16810_ = b[183:176];
      57'b?????????????????????????????????1???????????????????????:
        _16810_ = b[191:184];
      57'b????????????????????????????????1????????????????????????:
        _16810_ = b[199:192];
      57'b???????????????????????????????1?????????????????????????:
        _16810_ = b[207:200];
      57'b??????????????????????????????1??????????????????????????:
        _16810_ = b[215:208];
      57'b?????????????????????????????1???????????????????????????:
        _16810_ = b[223:216];
      57'b????????????????????????????1????????????????????????????:
        _16810_ = b[231:224];
      57'b???????????????????????????1?????????????????????????????:
        _16810_ = b[239:232];
      57'b??????????????????????????1??????????????????????????????:
        _16810_ = b[247:240];
      57'b?????????????????????????1???????????????????????????????:
        _16810_ = b[255:248];
      57'b????????????????????????1????????????????????????????????:
        _16810_ = b[263:256];
      57'b???????????????????????1?????????????????????????????????:
        _16810_ = b[271:264];
      57'b??????????????????????1??????????????????????????????????:
        _16810_ = b[279:272];
      57'b?????????????????????1???????????????????????????????????:
        _16810_ = b[287:280];
      57'b????????????????????1????????????????????????????????????:
        _16810_ = b[295:288];
      57'b???????????????????1?????????????????????????????????????:
        _16810_ = b[303:296];
      57'b??????????????????1??????????????????????????????????????:
        _16810_ = b[311:304];
      57'b?????????????????1???????????????????????????????????????:
        _16810_ = b[319:312];
      57'b????????????????1????????????????????????????????????????:
        _16810_ = b[327:320];
      57'b???????????????1?????????????????????????????????????????:
        _16810_ = b[335:328];
      57'b??????????????1??????????????????????????????????????????:
        _16810_ = b[343:336];
      57'b?????????????1???????????????????????????????????????????:
        _16810_ = b[351:344];
      57'b????????????1????????????????????????????????????????????:
        _16810_ = b[359:352];
      57'b???????????1?????????????????????????????????????????????:
        _16810_ = b[367:360];
      57'b??????????1??????????????????????????????????????????????:
        _16810_ = b[375:368];
      57'b?????????1???????????????????????????????????????????????:
        _16810_ = b[383:376];
      57'b????????1????????????????????????????????????????????????:
        _16810_ = b[391:384];
      57'b???????1?????????????????????????????????????????????????:
        _16810_ = b[399:392];
      57'b??????1??????????????????????????????????????????????????:
        _16810_ = b[407:400];
      57'b?????1???????????????????????????????????????????????????:
        _16810_ = b[415:408];
      57'b????1????????????????????????????????????????????????????:
        _16810_ = b[423:416];
      57'b???1?????????????????????????????????????????????????????:
        _16810_ = b[431:424];
      57'b??1??????????????????????????????????????????????????????:
        _16810_ = b[439:432];
      57'b?1???????????????????????????????????????????????????????:
        _16810_ = b[447:440];
      57'b1????????????????????????????????????????????????????????:
        _16810_ = b[455:448];
      default:
        _16810_ = a;
    endcase
  endfunction
  assign vec_data_056 = _16810_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440], data_d1[455:448] }, { _07405_, _07404_, _07403_, _07402_, _07401_, _07400_, _07399_, _07398_, _07397_, _07396_, _07395_, _07394_, _07393_, _07392_, _07391_, _07390_, _07389_, _07388_, _07387_, _07386_, _07385_, _07384_, _07383_, _07382_, _07381_, _07380_, _07379_, _07378_, _07377_, _07376_, _07375_, _07374_, _07373_, _07372_, _07371_, _07370_, _07369_, _07368_, _07367_, _07366_, _07365_, _07364_, _07363_, _07362_, _07361_, _07360_, _07359_, _07358_, _07357_, _07356_, _07355_, _07354_, _07353_, _07352_, _07351_, _07350_, _07349_ });
  assign _07349_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b111001;
  assign _07350_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b111000;
  assign _07351_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110111;
  assign _07352_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110110;
  assign _07353_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110101;
  assign _07354_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110100;
  assign _07355_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110011;
  assign _07356_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110010;
  assign _07357_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110001;
  assign _07358_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b110000;
  assign _07359_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101111;
  assign _07360_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101110;
  assign _07361_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101101;
  assign _07362_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101100;
  assign _07363_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101011;
  assign _07364_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101010;
  assign _07365_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101001;
  assign _07366_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b101000;
  assign _07367_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100111;
  assign _07368_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100110;
  assign _07369_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100101;
  assign _07370_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100100;
  assign _07371_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100011;
  assign _07372_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100010;
  assign _07373_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100001;
  assign _07374_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 6'b100000;
  assign _07375_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11111;
  assign _07376_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11110;
  assign _07377_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11101;
  assign _07378_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11100;
  assign _07379_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11011;
  assign _07380_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11010;
  assign _07381_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11001;
  assign _07382_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b11000;
  assign _07383_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10111;
  assign _07384_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10110;
  assign _07385_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10101;
  assign _07386_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10100;
  assign _07387_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10011;
  assign _07388_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10010;
  assign _07389_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10001;
  assign _07390_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 5'b10000;
  assign _07391_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1111;
  assign _07392_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1110;
  assign _07393_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1101;
  assign _07394_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1100;
  assign _07395_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1011;
  assign _07396_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1010;
  assign _07397_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1001;
  assign _07398_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 4'b1000;
  assign _07399_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 3'b111;
  assign _07400_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 3'b110;
  assign _07401_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 3'b101;
  assign _07402_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 3'b100;
  assign _07403_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 2'b11;
  assign _07404_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 2'b10;
  assign _07405_ = vec_sum_056_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5935" *) 1'b1;
  function [7:0] _16868_;
    input [7:0] a;
    input [447:0] b;
    input [55:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *)
    (* parallel_case *)
    casez (s)
      56'b???????????????????????????????????????????????????????1:
        _16868_ = b[7:0];
      56'b??????????????????????????????????????????????????????1?:
        _16868_ = b[15:8];
      56'b?????????????????????????????????????????????????????1??:
        _16868_ = b[23:16];
      56'b????????????????????????????????????????????????????1???:
        _16868_ = b[31:24];
      56'b???????????????????????????????????????????????????1????:
        _16868_ = b[39:32];
      56'b??????????????????????????????????????????????????1?????:
        _16868_ = b[47:40];
      56'b?????????????????????????????????????????????????1??????:
        _16868_ = b[55:48];
      56'b????????????????????????????????????????????????1???????:
        _16868_ = b[63:56];
      56'b???????????????????????????????????????????????1????????:
        _16868_ = b[71:64];
      56'b??????????????????????????????????????????????1?????????:
        _16868_ = b[79:72];
      56'b?????????????????????????????????????????????1??????????:
        _16868_ = b[87:80];
      56'b????????????????????????????????????????????1???????????:
        _16868_ = b[95:88];
      56'b???????????????????????????????????????????1????????????:
        _16868_ = b[103:96];
      56'b??????????????????????????????????????????1?????????????:
        _16868_ = b[111:104];
      56'b?????????????????????????????????????????1??????????????:
        _16868_ = b[119:112];
      56'b????????????????????????????????????????1???????????????:
        _16868_ = b[127:120];
      56'b???????????????????????????????????????1????????????????:
        _16868_ = b[135:128];
      56'b??????????????????????????????????????1?????????????????:
        _16868_ = b[143:136];
      56'b?????????????????????????????????????1??????????????????:
        _16868_ = b[151:144];
      56'b????????????????????????????????????1???????????????????:
        _16868_ = b[159:152];
      56'b???????????????????????????????????1????????????????????:
        _16868_ = b[167:160];
      56'b??????????????????????????????????1?????????????????????:
        _16868_ = b[175:168];
      56'b?????????????????????????????????1??????????????????????:
        _16868_ = b[183:176];
      56'b????????????????????????????????1???????????????????????:
        _16868_ = b[191:184];
      56'b???????????????????????????????1????????????????????????:
        _16868_ = b[199:192];
      56'b??????????????????????????????1?????????????????????????:
        _16868_ = b[207:200];
      56'b?????????????????????????????1??????????????????????????:
        _16868_ = b[215:208];
      56'b????????????????????????????1???????????????????????????:
        _16868_ = b[223:216];
      56'b???????????????????????????1????????????????????????????:
        _16868_ = b[231:224];
      56'b??????????????????????????1?????????????????????????????:
        _16868_ = b[239:232];
      56'b?????????????????????????1??????????????????????????????:
        _16868_ = b[247:240];
      56'b????????????????????????1???????????????????????????????:
        _16868_ = b[255:248];
      56'b???????????????????????1????????????????????????????????:
        _16868_ = b[263:256];
      56'b??????????????????????1?????????????????????????????????:
        _16868_ = b[271:264];
      56'b?????????????????????1??????????????????????????????????:
        _16868_ = b[279:272];
      56'b????????????????????1???????????????????????????????????:
        _16868_ = b[287:280];
      56'b???????????????????1????????????????????????????????????:
        _16868_ = b[295:288];
      56'b??????????????????1?????????????????????????????????????:
        _16868_ = b[303:296];
      56'b?????????????????1??????????????????????????????????????:
        _16868_ = b[311:304];
      56'b????????????????1???????????????????????????????????????:
        _16868_ = b[319:312];
      56'b???????????????1????????????????????????????????????????:
        _16868_ = b[327:320];
      56'b??????????????1?????????????????????????????????????????:
        _16868_ = b[335:328];
      56'b?????????????1??????????????????????????????????????????:
        _16868_ = b[343:336];
      56'b????????????1???????????????????????????????????????????:
        _16868_ = b[351:344];
      56'b???????????1????????????????????????????????????????????:
        _16868_ = b[359:352];
      56'b??????????1?????????????????????????????????????????????:
        _16868_ = b[367:360];
      56'b?????????1??????????????????????????????????????????????:
        _16868_ = b[375:368];
      56'b????????1???????????????????????????????????????????????:
        _16868_ = b[383:376];
      56'b???????1????????????????????????????????????????????????:
        _16868_ = b[391:384];
      56'b??????1?????????????????????????????????????????????????:
        _16868_ = b[399:392];
      56'b?????1??????????????????????????????????????????????????:
        _16868_ = b[407:400];
      56'b????1???????????????????????????????????????????????????:
        _16868_ = b[415:408];
      56'b???1????????????????????????????????????????????????????:
        _16868_ = b[423:416];
      56'b??1?????????????????????????????????????????????????????:
        _16868_ = b[431:424];
      56'b?1??????????????????????????????????????????????????????:
        _16868_ = b[439:432];
      56'b1???????????????????????????????????????????????????????:
        _16868_ = b[447:440];
      default:
        _16868_ = a;
    endcase
  endfunction
  assign vec_data_055 = _16868_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432], data_d1[447:440] }, { _07461_, _07460_, _07459_, _07458_, _07457_, _07456_, _07455_, _07454_, _07453_, _07452_, _07451_, _07450_, _07449_, _07448_, _07447_, _07446_, _07445_, _07444_, _07443_, _07442_, _07441_, _07440_, _07439_, _07438_, _07437_, _07436_, _07435_, _07434_, _07433_, _07432_, _07431_, _07430_, _07429_, _07428_, _07427_, _07426_, _07425_, _07424_, _07423_, _07422_, _07421_, _07420_, _07419_, _07418_, _07417_, _07416_, _07415_, _07414_, _07413_, _07412_, _07411_, _07410_, _07409_, _07408_, _07407_, _07406_ });
  assign _07406_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b111000;
  assign _07407_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110111;
  assign _07408_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110110;
  assign _07409_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110101;
  assign _07410_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110100;
  assign _07411_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110011;
  assign _07412_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110010;
  assign _07413_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110001;
  assign _07414_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b110000;
  assign _07415_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101111;
  assign _07416_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101110;
  assign _07417_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101101;
  assign _07418_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101100;
  assign _07419_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101011;
  assign _07420_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101010;
  assign _07421_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101001;
  assign _07422_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b101000;
  assign _07423_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100111;
  assign _07424_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100110;
  assign _07425_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100101;
  assign _07426_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100100;
  assign _07427_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100011;
  assign _07428_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100010;
  assign _07429_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100001;
  assign _07430_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 6'b100000;
  assign _07431_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11111;
  assign _07432_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11110;
  assign _07433_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11101;
  assign _07434_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11100;
  assign _07435_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11011;
  assign _07436_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11010;
  assign _07437_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11001;
  assign _07438_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b11000;
  assign _07439_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10111;
  assign _07440_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10110;
  assign _07441_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10101;
  assign _07442_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10100;
  assign _07443_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5890|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10011;
  assign _07444_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5889|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10010;
  assign _07445_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5888|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10001;
  assign _07446_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5887|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 5'b10000;
  assign _07447_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5886|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1111;
  assign _07448_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5885|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1110;
  assign _07449_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5884|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1101;
  assign _07450_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5883|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1100;
  assign _07451_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1011;
  assign _07452_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1010;
  assign _07453_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1001;
  assign _07454_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 4'b1000;
  assign _07455_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 3'b111;
  assign _07456_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 3'b110;
  assign _07457_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 3'b101;
  assign _07458_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 3'b100;
  assign _07459_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 2'b11;
  assign _07460_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 2'b10;
  assign _07461_ = vec_sum_055_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5871" *) 1'b1;
  function [7:0] _16925_;
    input [7:0] a;
    input [439:0] b;
    input [54:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *)
    (* parallel_case *)
    casez (s)
      55'b??????????????????????????????????????????????????????1:
        _16925_ = b[7:0];
      55'b?????????????????????????????????????????????????????1?:
        _16925_ = b[15:8];
      55'b????????????????????????????????????????????????????1??:
        _16925_ = b[23:16];
      55'b???????????????????????????????????????????????????1???:
        _16925_ = b[31:24];
      55'b??????????????????????????????????????????????????1????:
        _16925_ = b[39:32];
      55'b?????????????????????????????????????????????????1?????:
        _16925_ = b[47:40];
      55'b????????????????????????????????????????????????1??????:
        _16925_ = b[55:48];
      55'b???????????????????????????????????????????????1???????:
        _16925_ = b[63:56];
      55'b??????????????????????????????????????????????1????????:
        _16925_ = b[71:64];
      55'b?????????????????????????????????????????????1?????????:
        _16925_ = b[79:72];
      55'b????????????????????????????????????????????1??????????:
        _16925_ = b[87:80];
      55'b???????????????????????????????????????????1???????????:
        _16925_ = b[95:88];
      55'b??????????????????????????????????????????1????????????:
        _16925_ = b[103:96];
      55'b?????????????????????????????????????????1?????????????:
        _16925_ = b[111:104];
      55'b????????????????????????????????????????1??????????????:
        _16925_ = b[119:112];
      55'b???????????????????????????????????????1???????????????:
        _16925_ = b[127:120];
      55'b??????????????????????????????????????1????????????????:
        _16925_ = b[135:128];
      55'b?????????????????????????????????????1?????????????????:
        _16925_ = b[143:136];
      55'b????????????????????????????????????1??????????????????:
        _16925_ = b[151:144];
      55'b???????????????????????????????????1???????????????????:
        _16925_ = b[159:152];
      55'b??????????????????????????????????1????????????????????:
        _16925_ = b[167:160];
      55'b?????????????????????????????????1?????????????????????:
        _16925_ = b[175:168];
      55'b????????????????????????????????1??????????????????????:
        _16925_ = b[183:176];
      55'b???????????????????????????????1???????????????????????:
        _16925_ = b[191:184];
      55'b??????????????????????????????1????????????????????????:
        _16925_ = b[199:192];
      55'b?????????????????????????????1?????????????????????????:
        _16925_ = b[207:200];
      55'b????????????????????????????1??????????????????????????:
        _16925_ = b[215:208];
      55'b???????????????????????????1???????????????????????????:
        _16925_ = b[223:216];
      55'b??????????????????????????1????????????????????????????:
        _16925_ = b[231:224];
      55'b?????????????????????????1?????????????????????????????:
        _16925_ = b[239:232];
      55'b????????????????????????1??????????????????????????????:
        _16925_ = b[247:240];
      55'b???????????????????????1???????????????????????????????:
        _16925_ = b[255:248];
      55'b??????????????????????1????????????????????????????????:
        _16925_ = b[263:256];
      55'b?????????????????????1?????????????????????????????????:
        _16925_ = b[271:264];
      55'b????????????????????1??????????????????????????????????:
        _16925_ = b[279:272];
      55'b???????????????????1???????????????????????????????????:
        _16925_ = b[287:280];
      55'b??????????????????1????????????????????????????????????:
        _16925_ = b[295:288];
      55'b?????????????????1?????????????????????????????????????:
        _16925_ = b[303:296];
      55'b????????????????1??????????????????????????????????????:
        _16925_ = b[311:304];
      55'b???????????????1???????????????????????????????????????:
        _16925_ = b[319:312];
      55'b??????????????1????????????????????????????????????????:
        _16925_ = b[327:320];
      55'b?????????????1?????????????????????????????????????????:
        _16925_ = b[335:328];
      55'b????????????1??????????????????????????????????????????:
        _16925_ = b[343:336];
      55'b???????????1???????????????????????????????????????????:
        _16925_ = b[351:344];
      55'b??????????1????????????????????????????????????????????:
        _16925_ = b[359:352];
      55'b?????????1?????????????????????????????????????????????:
        _16925_ = b[367:360];
      55'b????????1??????????????????????????????????????????????:
        _16925_ = b[375:368];
      55'b???????1???????????????????????????????????????????????:
        _16925_ = b[383:376];
      55'b??????1????????????????????????????????????????????????:
        _16925_ = b[391:384];
      55'b?????1?????????????????????????????????????????????????:
        _16925_ = b[399:392];
      55'b????1??????????????????????????????????????????????????:
        _16925_ = b[407:400];
      55'b???1???????????????????????????????????????????????????:
        _16925_ = b[415:408];
      55'b??1????????????????????????????????????????????????????:
        _16925_ = b[423:416];
      55'b?1?????????????????????????????????????????????????????:
        _16925_ = b[431:424];
      55'b1??????????????????????????????????????????????????????:
        _16925_ = b[439:432];
      default:
        _16925_ = a;
    endcase
  endfunction
  assign vec_data_054 = _16925_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424], data_d1[439:432] }, { _07516_, _07515_, _07514_, _07513_, _07512_, _07511_, _07510_, _07509_, _07508_, _07507_, _07506_, _07505_, _07504_, _07503_, _07502_, _07501_, _07500_, _07499_, _07498_, _07497_, _07496_, _07495_, _07494_, _07493_, _07492_, _07491_, _07490_, _07489_, _07488_, _07487_, _07486_, _07485_, _07484_, _07483_, _07482_, _07481_, _07480_, _07479_, _07478_, _07477_, _07476_, _07475_, _07474_, _07473_, _07472_, _07471_, _07470_, _07469_, _07468_, _07467_, _07466_, _07465_, _07464_, _07463_, _07462_ });
  assign _07462_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110111;
  assign _07463_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110110;
  assign _07464_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110101;
  assign _07465_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110100;
  assign _07466_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110011;
  assign _07467_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110010;
  assign _07468_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110001;
  assign _07469_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b110000;
  assign _07470_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101111;
  assign _07471_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101110;
  assign _07472_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101101;
  assign _07473_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101100;
  assign _07474_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101011;
  assign _07475_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101010;
  assign _07476_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101001;
  assign _07477_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b101000;
  assign _07478_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100111;
  assign _07479_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100110;
  assign _07480_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5845|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100101;
  assign _07481_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5844|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100100;
  assign _07482_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5843|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100011;
  assign _07483_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5842|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100010;
  assign _07484_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5841|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100001;
  assign _07485_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5840|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 6'b100000;
  assign _07486_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5839|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11111;
  assign _07487_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5838|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11110;
  assign _07488_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11101;
  assign _07489_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11100;
  assign _07490_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11011;
  assign _07491_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11010;
  assign _07492_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11001;
  assign _07493_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b11000;
  assign _07494_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10111;
  assign _07495_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10110;
  assign _07496_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10101;
  assign _07497_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10100;
  assign _07498_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10011;
  assign _07499_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10010;
  assign _07500_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10001;
  assign _07501_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 5'b10000;
  assign _07502_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1111;
  assign _07503_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1110;
  assign _07504_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1101;
  assign _07505_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1100;
  assign _07506_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1011;
  assign _07507_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1010;
  assign _07508_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1001;
  assign _07509_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 4'b1000;
  assign _07510_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 3'b111;
  assign _07511_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 3'b110;
  assign _07512_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 3'b101;
  assign _07513_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 3'b100;
  assign _07514_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 2'b11;
  assign _07515_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 2'b10;
  assign _07516_ = vec_sum_054_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5808" *) 1'b1;
  function [7:0] _16981_;
    input [7:0] a;
    input [431:0] b;
    input [53:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *)
    (* parallel_case *)
    casez (s)
      54'b?????????????????????????????????????????????????????1:
        _16981_ = b[7:0];
      54'b????????????????????????????????????????????????????1?:
        _16981_ = b[15:8];
      54'b???????????????????????????????????????????????????1??:
        _16981_ = b[23:16];
      54'b??????????????????????????????????????????????????1???:
        _16981_ = b[31:24];
      54'b?????????????????????????????????????????????????1????:
        _16981_ = b[39:32];
      54'b????????????????????????????????????????????????1?????:
        _16981_ = b[47:40];
      54'b???????????????????????????????????????????????1??????:
        _16981_ = b[55:48];
      54'b??????????????????????????????????????????????1???????:
        _16981_ = b[63:56];
      54'b?????????????????????????????????????????????1????????:
        _16981_ = b[71:64];
      54'b????????????????????????????????????????????1?????????:
        _16981_ = b[79:72];
      54'b???????????????????????????????????????????1??????????:
        _16981_ = b[87:80];
      54'b??????????????????????????????????????????1???????????:
        _16981_ = b[95:88];
      54'b?????????????????????????????????????????1????????????:
        _16981_ = b[103:96];
      54'b????????????????????????????????????????1?????????????:
        _16981_ = b[111:104];
      54'b???????????????????????????????????????1??????????????:
        _16981_ = b[119:112];
      54'b??????????????????????????????????????1???????????????:
        _16981_ = b[127:120];
      54'b?????????????????????????????????????1????????????????:
        _16981_ = b[135:128];
      54'b????????????????????????????????????1?????????????????:
        _16981_ = b[143:136];
      54'b???????????????????????????????????1??????????????????:
        _16981_ = b[151:144];
      54'b??????????????????????????????????1???????????????????:
        _16981_ = b[159:152];
      54'b?????????????????????????????????1????????????????????:
        _16981_ = b[167:160];
      54'b????????????????????????????????1?????????????????????:
        _16981_ = b[175:168];
      54'b???????????????????????????????1??????????????????????:
        _16981_ = b[183:176];
      54'b??????????????????????????????1???????????????????????:
        _16981_ = b[191:184];
      54'b?????????????????????????????1????????????????????????:
        _16981_ = b[199:192];
      54'b????????????????????????????1?????????????????????????:
        _16981_ = b[207:200];
      54'b???????????????????????????1??????????????????????????:
        _16981_ = b[215:208];
      54'b??????????????????????????1???????????????????????????:
        _16981_ = b[223:216];
      54'b?????????????????????????1????????????????????????????:
        _16981_ = b[231:224];
      54'b????????????????????????1?????????????????????????????:
        _16981_ = b[239:232];
      54'b???????????????????????1??????????????????????????????:
        _16981_ = b[247:240];
      54'b??????????????????????1???????????????????????????????:
        _16981_ = b[255:248];
      54'b?????????????????????1????????????????????????????????:
        _16981_ = b[263:256];
      54'b????????????????????1?????????????????????????????????:
        _16981_ = b[271:264];
      54'b???????????????????1??????????????????????????????????:
        _16981_ = b[279:272];
      54'b??????????????????1???????????????????????????????????:
        _16981_ = b[287:280];
      54'b?????????????????1????????????????????????????????????:
        _16981_ = b[295:288];
      54'b????????????????1?????????????????????????????????????:
        _16981_ = b[303:296];
      54'b???????????????1??????????????????????????????????????:
        _16981_ = b[311:304];
      54'b??????????????1???????????????????????????????????????:
        _16981_ = b[319:312];
      54'b?????????????1????????????????????????????????????????:
        _16981_ = b[327:320];
      54'b????????????1?????????????????????????????????????????:
        _16981_ = b[335:328];
      54'b???????????1??????????????????????????????????????????:
        _16981_ = b[343:336];
      54'b??????????1???????????????????????????????????????????:
        _16981_ = b[351:344];
      54'b?????????1????????????????????????????????????????????:
        _16981_ = b[359:352];
      54'b????????1?????????????????????????????????????????????:
        _16981_ = b[367:360];
      54'b???????1??????????????????????????????????????????????:
        _16981_ = b[375:368];
      54'b??????1???????????????????????????????????????????????:
        _16981_ = b[383:376];
      54'b?????1????????????????????????????????????????????????:
        _16981_ = b[391:384];
      54'b????1?????????????????????????????????????????????????:
        _16981_ = b[399:392];
      54'b???1??????????????????????????????????????????????????:
        _16981_ = b[407:400];
      54'b??1???????????????????????????????????????????????????:
        _16981_ = b[415:408];
      54'b?1????????????????????????????????????????????????????:
        _16981_ = b[423:416];
      54'b1?????????????????????????????????????????????????????:
        _16981_ = b[431:424];
      default:
        _16981_ = a;
    endcase
  endfunction
  assign vec_data_053 = _16981_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416], data_d1[431:424] }, { _07570_, _07569_, _07568_, _07567_, _07566_, _07565_, _07564_, _07563_, _07562_, _07561_, _07560_, _07559_, _07558_, _07557_, _07556_, _07555_, _07554_, _07553_, _07552_, _07551_, _07550_, _07549_, _07548_, _07547_, _07546_, _07545_, _07544_, _07543_, _07542_, _07541_, _07540_, _07539_, _07538_, _07537_, _07536_, _07535_, _07534_, _07533_, _07532_, _07531_, _07530_, _07529_, _07528_, _07527_, _07526_, _07525_, _07524_, _07523_, _07522_, _07521_, _07520_, _07519_, _07518_, _07517_ });
  assign _07517_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5800|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110110;
  assign _07518_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5799|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110101;
  assign _07519_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5798|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110100;
  assign _07520_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5797|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110011;
  assign _07521_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5796|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110010;
  assign _07522_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5795|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110001;
  assign _07523_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5794|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b110000;
  assign _07524_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101111;
  assign _07525_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101110;
  assign _07526_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101101;
  assign _07527_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101100;
  assign _07528_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101011;
  assign _07529_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101010;
  assign _07530_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101001;
  assign _07531_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b101000;
  assign _07532_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100111;
  assign _07533_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100110;
  assign _07534_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100101;
  assign _07535_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100100;
  assign _07536_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100011;
  assign _07537_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100010;
  assign _07538_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100001;
  assign _07539_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 6'b100000;
  assign _07540_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11111;
  assign _07541_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11110;
  assign _07542_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11101;
  assign _07543_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11100;
  assign _07544_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11011;
  assign _07545_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11010;
  assign _07546_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11001;
  assign _07547_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b11000;
  assign _07548_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10111;
  assign _07549_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10110;
  assign _07550_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10101;
  assign _07551_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10100;
  assign _07552_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10011;
  assign _07553_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10010;
  assign _07554_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10001;
  assign _07555_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 5'b10000;
  assign _07556_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1111;
  assign _07557_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1110;
  assign _07558_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1101;
  assign _07559_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5758|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1100;
  assign _07560_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5757|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1011;
  assign _07561_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5756|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1010;
  assign _07562_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5755|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1001;
  assign _07563_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5754|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 4'b1000;
  assign _07564_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5753|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 3'b111;
  assign _07565_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5752|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 3'b110;
  assign _07566_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5751|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 3'b101;
  assign _07567_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 3'b100;
  assign _07568_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 2'b11;
  assign _07569_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 2'b10;
  assign _07570_ = vec_sum_053_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5746" *) 1'b1;
  function [7:0] _17036_;
    input [7:0] a;
    input [423:0] b;
    input [52:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *)
    (* parallel_case *)
    casez (s)
      53'b????????????????????????????????????????????????????1:
        _17036_ = b[7:0];
      53'b???????????????????????????????????????????????????1?:
        _17036_ = b[15:8];
      53'b??????????????????????????????????????????????????1??:
        _17036_ = b[23:16];
      53'b?????????????????????????????????????????????????1???:
        _17036_ = b[31:24];
      53'b????????????????????????????????????????????????1????:
        _17036_ = b[39:32];
      53'b???????????????????????????????????????????????1?????:
        _17036_ = b[47:40];
      53'b??????????????????????????????????????????????1??????:
        _17036_ = b[55:48];
      53'b?????????????????????????????????????????????1???????:
        _17036_ = b[63:56];
      53'b????????????????????????????????????????????1????????:
        _17036_ = b[71:64];
      53'b???????????????????????????????????????????1?????????:
        _17036_ = b[79:72];
      53'b??????????????????????????????????????????1??????????:
        _17036_ = b[87:80];
      53'b?????????????????????????????????????????1???????????:
        _17036_ = b[95:88];
      53'b????????????????????????????????????????1????????????:
        _17036_ = b[103:96];
      53'b???????????????????????????????????????1?????????????:
        _17036_ = b[111:104];
      53'b??????????????????????????????????????1??????????????:
        _17036_ = b[119:112];
      53'b?????????????????????????????????????1???????????????:
        _17036_ = b[127:120];
      53'b????????????????????????????????????1????????????????:
        _17036_ = b[135:128];
      53'b???????????????????????????????????1?????????????????:
        _17036_ = b[143:136];
      53'b??????????????????????????????????1??????????????????:
        _17036_ = b[151:144];
      53'b?????????????????????????????????1???????????????????:
        _17036_ = b[159:152];
      53'b????????????????????????????????1????????????????????:
        _17036_ = b[167:160];
      53'b???????????????????????????????1?????????????????????:
        _17036_ = b[175:168];
      53'b??????????????????????????????1??????????????????????:
        _17036_ = b[183:176];
      53'b?????????????????????????????1???????????????????????:
        _17036_ = b[191:184];
      53'b????????????????????????????1????????????????????????:
        _17036_ = b[199:192];
      53'b???????????????????????????1?????????????????????????:
        _17036_ = b[207:200];
      53'b??????????????????????????1??????????????????????????:
        _17036_ = b[215:208];
      53'b?????????????????????????1???????????????????????????:
        _17036_ = b[223:216];
      53'b????????????????????????1????????????????????????????:
        _17036_ = b[231:224];
      53'b???????????????????????1?????????????????????????????:
        _17036_ = b[239:232];
      53'b??????????????????????1??????????????????????????????:
        _17036_ = b[247:240];
      53'b?????????????????????1???????????????????????????????:
        _17036_ = b[255:248];
      53'b????????????????????1????????????????????????????????:
        _17036_ = b[263:256];
      53'b???????????????????1?????????????????????????????????:
        _17036_ = b[271:264];
      53'b??????????????????1??????????????????????????????????:
        _17036_ = b[279:272];
      53'b?????????????????1???????????????????????????????????:
        _17036_ = b[287:280];
      53'b????????????????1????????????????????????????????????:
        _17036_ = b[295:288];
      53'b???????????????1?????????????????????????????????????:
        _17036_ = b[303:296];
      53'b??????????????1??????????????????????????????????????:
        _17036_ = b[311:304];
      53'b?????????????1???????????????????????????????????????:
        _17036_ = b[319:312];
      53'b????????????1????????????????????????????????????????:
        _17036_ = b[327:320];
      53'b???????????1?????????????????????????????????????????:
        _17036_ = b[335:328];
      53'b??????????1??????????????????????????????????????????:
        _17036_ = b[343:336];
      53'b?????????1???????????????????????????????????????????:
        _17036_ = b[351:344];
      53'b????????1????????????????????????????????????????????:
        _17036_ = b[359:352];
      53'b???????1?????????????????????????????????????????????:
        _17036_ = b[367:360];
      53'b??????1??????????????????????????????????????????????:
        _17036_ = b[375:368];
      53'b?????1???????????????????????????????????????????????:
        _17036_ = b[383:376];
      53'b????1????????????????????????????????????????????????:
        _17036_ = b[391:384];
      53'b???1?????????????????????????????????????????????????:
        _17036_ = b[399:392];
      53'b??1??????????????????????????????????????????????????:
        _17036_ = b[407:400];
      53'b?1???????????????????????????????????????????????????:
        _17036_ = b[415:408];
      53'b1????????????????????????????????????????????????????:
        _17036_ = b[423:416];
      default:
        _17036_ = a;
    endcase
  endfunction
  assign vec_data_052 = _17036_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408], data_d1[423:416] }, { _07623_, _07622_, _07621_, _07620_, _07619_, _07618_, _07617_, _07616_, _07615_, _07614_, _07613_, _07612_, _07611_, _07610_, _07609_, _07608_, _07607_, _07606_, _07605_, _07604_, _07603_, _07602_, _07601_, _07600_, _07599_, _07598_, _07597_, _07596_, _07595_, _07594_, _07593_, _07592_, _07591_, _07590_, _07589_, _07588_, _07587_, _07586_, _07585_, _07584_, _07583_, _07582_, _07581_, _07580_, _07579_, _07578_, _07577_, _07576_, _07575_, _07574_, _07573_, _07572_, _07571_ });
  assign _07571_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110101;
  assign _07572_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110100;
  assign _07573_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110011;
  assign _07574_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110010;
  assign _07575_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110001;
  assign _07576_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b110000;
  assign _07577_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101111;
  assign _07578_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101110;
  assign _07579_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101101;
  assign _07580_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101100;
  assign _07581_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101011;
  assign _07582_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101010;
  assign _07583_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101001;
  assign _07584_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b101000;
  assign _07585_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100111;
  assign _07586_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100110;
  assign _07587_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100101;
  assign _07588_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100100;
  assign _07589_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100011;
  assign _07590_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100010;
  assign _07591_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100001;
  assign _07592_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 6'b100000;
  assign _07593_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5716|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11111;
  assign _07594_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5715|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11110;
  assign _07595_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5714|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11101;
  assign _07596_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5713|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11100;
  assign _07597_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5712|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11011;
  assign _07598_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5711|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11010;
  assign _07599_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5710|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11001;
  assign _07600_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5709|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b11000;
  assign _07601_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10111;
  assign _07602_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10110;
  assign _07603_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10101;
  assign _07604_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10100;
  assign _07605_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10011;
  assign _07606_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10010;
  assign _07607_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10001;
  assign _07608_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 5'b10000;
  assign _07609_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1111;
  assign _07610_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1110;
  assign _07611_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1101;
  assign _07612_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1100;
  assign _07613_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1011;
  assign _07614_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1010;
  assign _07615_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1001;
  assign _07616_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 4'b1000;
  assign _07617_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 3'b111;
  assign _07618_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 3'b110;
  assign _07619_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 3'b101;
  assign _07620_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 3'b100;
  assign _07621_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 2'b11;
  assign _07622_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 2'b10;
  assign _07623_ = vec_sum_052_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5685" *) 1'b1;
  function [7:0] _17090_;
    input [7:0] a;
    input [415:0] b;
    input [51:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *)
    (* parallel_case *)
    casez (s)
      52'b???????????????????????????????????????????????????1:
        _17090_ = b[7:0];
      52'b??????????????????????????????????????????????????1?:
        _17090_ = b[15:8];
      52'b?????????????????????????????????????????????????1??:
        _17090_ = b[23:16];
      52'b????????????????????????????????????????????????1???:
        _17090_ = b[31:24];
      52'b???????????????????????????????????????????????1????:
        _17090_ = b[39:32];
      52'b??????????????????????????????????????????????1?????:
        _17090_ = b[47:40];
      52'b?????????????????????????????????????????????1??????:
        _17090_ = b[55:48];
      52'b????????????????????????????????????????????1???????:
        _17090_ = b[63:56];
      52'b???????????????????????????????????????????1????????:
        _17090_ = b[71:64];
      52'b??????????????????????????????????????????1?????????:
        _17090_ = b[79:72];
      52'b?????????????????????????????????????????1??????????:
        _17090_ = b[87:80];
      52'b????????????????????????????????????????1???????????:
        _17090_ = b[95:88];
      52'b???????????????????????????????????????1????????????:
        _17090_ = b[103:96];
      52'b??????????????????????????????????????1?????????????:
        _17090_ = b[111:104];
      52'b?????????????????????????????????????1??????????????:
        _17090_ = b[119:112];
      52'b????????????????????????????????????1???????????????:
        _17090_ = b[127:120];
      52'b???????????????????????????????????1????????????????:
        _17090_ = b[135:128];
      52'b??????????????????????????????????1?????????????????:
        _17090_ = b[143:136];
      52'b?????????????????????????????????1??????????????????:
        _17090_ = b[151:144];
      52'b????????????????????????????????1???????????????????:
        _17090_ = b[159:152];
      52'b???????????????????????????????1????????????????????:
        _17090_ = b[167:160];
      52'b??????????????????????????????1?????????????????????:
        _17090_ = b[175:168];
      52'b?????????????????????????????1??????????????????????:
        _17090_ = b[183:176];
      52'b????????????????????????????1???????????????????????:
        _17090_ = b[191:184];
      52'b???????????????????????????1????????????????????????:
        _17090_ = b[199:192];
      52'b??????????????????????????1?????????????????????????:
        _17090_ = b[207:200];
      52'b?????????????????????????1??????????????????????????:
        _17090_ = b[215:208];
      52'b????????????????????????1???????????????????????????:
        _17090_ = b[223:216];
      52'b???????????????????????1????????????????????????????:
        _17090_ = b[231:224];
      52'b??????????????????????1?????????????????????????????:
        _17090_ = b[239:232];
      52'b?????????????????????1??????????????????????????????:
        _17090_ = b[247:240];
      52'b????????????????????1???????????????????????????????:
        _17090_ = b[255:248];
      52'b???????????????????1????????????????????????????????:
        _17090_ = b[263:256];
      52'b??????????????????1?????????????????????????????????:
        _17090_ = b[271:264];
      52'b?????????????????1??????????????????????????????????:
        _17090_ = b[279:272];
      52'b????????????????1???????????????????????????????????:
        _17090_ = b[287:280];
      52'b???????????????1????????????????????????????????????:
        _17090_ = b[295:288];
      52'b??????????????1?????????????????????????????????????:
        _17090_ = b[303:296];
      52'b?????????????1??????????????????????????????????????:
        _17090_ = b[311:304];
      52'b????????????1???????????????????????????????????????:
        _17090_ = b[319:312];
      52'b???????????1????????????????????????????????????????:
        _17090_ = b[327:320];
      52'b??????????1?????????????????????????????????????????:
        _17090_ = b[335:328];
      52'b?????????1??????????????????????????????????????????:
        _17090_ = b[343:336];
      52'b????????1???????????????????????????????????????????:
        _17090_ = b[351:344];
      52'b???????1????????????????????????????????????????????:
        _17090_ = b[359:352];
      52'b??????1?????????????????????????????????????????????:
        _17090_ = b[367:360];
      52'b?????1??????????????????????????????????????????????:
        _17090_ = b[375:368];
      52'b????1???????????????????????????????????????????????:
        _17090_ = b[383:376];
      52'b???1????????????????????????????????????????????????:
        _17090_ = b[391:384];
      52'b??1?????????????????????????????????????????????????:
        _17090_ = b[399:392];
      52'b?1??????????????????????????????????????????????????:
        _17090_ = b[407:400];
      52'b1???????????????????????????????????????????????????:
        _17090_ = b[415:408];
      default:
        _17090_ = a;
    endcase
  endfunction
  assign vec_data_051 = _17090_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400], data_d1[415:408] }, { _07675_, _07674_, _07673_, _07672_, _07671_, _07670_, _07669_, _07668_, _07667_, _07666_, _07665_, _07664_, _07663_, _07662_, _07661_, _07660_, _07659_, _07658_, _07657_, _07656_, _07655_, _07654_, _07653_, _07652_, _07651_, _07650_, _07649_, _07648_, _07647_, _07646_, _07645_, _07644_, _07643_, _07642_, _07641_, _07640_, _07639_, _07638_, _07637_, _07636_, _07635_, _07634_, _07633_, _07632_, _07631_, _07630_, _07629_, _07628_, _07627_, _07626_, _07625_, _07624_ });
  assign _07624_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b110100;
  assign _07625_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b110011;
  assign _07626_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5675|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b110010;
  assign _07627_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5674|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b110001;
  assign _07628_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5673|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b110000;
  assign _07629_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5672|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101111;
  assign _07630_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5671|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101110;
  assign _07631_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5670|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101101;
  assign _07632_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5669|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101100;
  assign _07633_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5668|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101011;
  assign _07634_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101010;
  assign _07635_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101001;
  assign _07636_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b101000;
  assign _07637_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100111;
  assign _07638_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100110;
  assign _07639_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100101;
  assign _07640_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100100;
  assign _07641_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100011;
  assign _07642_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100010;
  assign _07643_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100001;
  assign _07644_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 6'b100000;
  assign _07645_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11111;
  assign _07646_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11110;
  assign _07647_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11101;
  assign _07648_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11100;
  assign _07649_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11011;
  assign _07650_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11010;
  assign _07651_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11001;
  assign _07652_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b11000;
  assign _07653_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10111;
  assign _07654_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10110;
  assign _07655_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10101;
  assign _07656_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10100;
  assign _07657_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10011;
  assign _07658_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10010;
  assign _07659_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10001;
  assign _07660_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 5'b10000;
  assign _07661_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1111;
  assign _07662_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1110;
  assign _07663_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1101;
  assign _07664_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1100;
  assign _07665_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1011;
  assign _07666_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5635|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1010;
  assign _07667_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5634|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1001;
  assign _07668_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5633|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 4'b1000;
  assign _07669_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5632|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 3'b111;
  assign _07670_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5631|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 3'b110;
  assign _07671_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5630|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 3'b101;
  assign _07672_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5629|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 3'b100;
  assign _07673_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5628|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 2'b11;
  assign _07674_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 2'b10;
  assign _07675_ = vec_sum_051_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5625" *) 1'b1;
  function [7:0] _17143_;
    input [7:0] a;
    input [407:0] b;
    input [50:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *)
    (* parallel_case *)
    casez (s)
      51'b??????????????????????????????????????????????????1:
        _17143_ = b[7:0];
      51'b?????????????????????????????????????????????????1?:
        _17143_ = b[15:8];
      51'b????????????????????????????????????????????????1??:
        _17143_ = b[23:16];
      51'b???????????????????????????????????????????????1???:
        _17143_ = b[31:24];
      51'b??????????????????????????????????????????????1????:
        _17143_ = b[39:32];
      51'b?????????????????????????????????????????????1?????:
        _17143_ = b[47:40];
      51'b????????????????????????????????????????????1??????:
        _17143_ = b[55:48];
      51'b???????????????????????????????????????????1???????:
        _17143_ = b[63:56];
      51'b??????????????????????????????????????????1????????:
        _17143_ = b[71:64];
      51'b?????????????????????????????????????????1?????????:
        _17143_ = b[79:72];
      51'b????????????????????????????????????????1??????????:
        _17143_ = b[87:80];
      51'b???????????????????????????????????????1???????????:
        _17143_ = b[95:88];
      51'b??????????????????????????????????????1????????????:
        _17143_ = b[103:96];
      51'b?????????????????????????????????????1?????????????:
        _17143_ = b[111:104];
      51'b????????????????????????????????????1??????????????:
        _17143_ = b[119:112];
      51'b???????????????????????????????????1???????????????:
        _17143_ = b[127:120];
      51'b??????????????????????????????????1????????????????:
        _17143_ = b[135:128];
      51'b?????????????????????????????????1?????????????????:
        _17143_ = b[143:136];
      51'b????????????????????????????????1??????????????????:
        _17143_ = b[151:144];
      51'b???????????????????????????????1???????????????????:
        _17143_ = b[159:152];
      51'b??????????????????????????????1????????????????????:
        _17143_ = b[167:160];
      51'b?????????????????????????????1?????????????????????:
        _17143_ = b[175:168];
      51'b????????????????????????????1??????????????????????:
        _17143_ = b[183:176];
      51'b???????????????????????????1???????????????????????:
        _17143_ = b[191:184];
      51'b??????????????????????????1????????????????????????:
        _17143_ = b[199:192];
      51'b?????????????????????????1?????????????????????????:
        _17143_ = b[207:200];
      51'b????????????????????????1??????????????????????????:
        _17143_ = b[215:208];
      51'b???????????????????????1???????????????????????????:
        _17143_ = b[223:216];
      51'b??????????????????????1????????????????????????????:
        _17143_ = b[231:224];
      51'b?????????????????????1?????????????????????????????:
        _17143_ = b[239:232];
      51'b????????????????????1??????????????????????????????:
        _17143_ = b[247:240];
      51'b???????????????????1???????????????????????????????:
        _17143_ = b[255:248];
      51'b??????????????????1????????????????????????????????:
        _17143_ = b[263:256];
      51'b?????????????????1?????????????????????????????????:
        _17143_ = b[271:264];
      51'b????????????????1??????????????????????????????????:
        _17143_ = b[279:272];
      51'b???????????????1???????????????????????????????????:
        _17143_ = b[287:280];
      51'b??????????????1????????????????????????????????????:
        _17143_ = b[295:288];
      51'b?????????????1?????????????????????????????????????:
        _17143_ = b[303:296];
      51'b????????????1??????????????????????????????????????:
        _17143_ = b[311:304];
      51'b???????????1???????????????????????????????????????:
        _17143_ = b[319:312];
      51'b??????????1????????????????????????????????????????:
        _17143_ = b[327:320];
      51'b?????????1?????????????????????????????????????????:
        _17143_ = b[335:328];
      51'b????????1??????????????????????????????????????????:
        _17143_ = b[343:336];
      51'b???????1???????????????????????????????????????????:
        _17143_ = b[351:344];
      51'b??????1????????????????????????????????????????????:
        _17143_ = b[359:352];
      51'b?????1?????????????????????????????????????????????:
        _17143_ = b[367:360];
      51'b????1??????????????????????????????????????????????:
        _17143_ = b[375:368];
      51'b???1???????????????????????????????????????????????:
        _17143_ = b[383:376];
      51'b??1????????????????????????????????????????????????:
        _17143_ = b[391:384];
      51'b?1?????????????????????????????????????????????????:
        _17143_ = b[399:392];
      51'b1??????????????????????????????????????????????????:
        _17143_ = b[407:400];
      default:
        _17143_ = a;
    endcase
  endfunction
  assign vec_data_050 = _17143_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392], data_d1[407:400] }, { _07726_, _07725_, _07724_, _07723_, _07722_, _07721_, _07720_, _07719_, _07718_, _07717_, _07716_, _07715_, _07714_, _07713_, _07712_, _07711_, _07710_, _07709_, _07708_, _07707_, _07706_, _07705_, _07704_, _07703_, _07702_, _07701_, _07700_, _07699_, _07698_, _07697_, _07696_, _07695_, _07694_, _07693_, _07692_, _07691_, _07690_, _07689_, _07688_, _07687_, _07686_, _07685_, _07684_, _07683_, _07682_, _07681_, _07680_, _07679_, _07678_, _07677_, _07676_ });
  assign _07676_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b110011;
  assign _07677_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b110010;
  assign _07678_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b110001;
  assign _07679_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b110000;
  assign _07680_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101111;
  assign _07681_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101110;
  assign _07682_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101101;
  assign _07683_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101100;
  assign _07684_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101011;
  assign _07685_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101010;
  assign _07686_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101001;
  assign _07687_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b101000;
  assign _07688_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100111;
  assign _07689_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100110;
  assign _07690_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100101;
  assign _07691_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100100;
  assign _07692_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100011;
  assign _07693_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100010;
  assign _07694_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100001;
  assign _07695_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 6'b100000;
  assign _07696_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11111;
  assign _07697_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5596|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11110;
  assign _07698_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5595|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11101;
  assign _07699_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5594|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11100;
  assign _07700_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5593|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11011;
  assign _07701_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5592|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11010;
  assign _07702_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5591|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11001;
  assign _07703_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5590|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b11000;
  assign _07704_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5589|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10111;
  assign _07705_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10110;
  assign _07706_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10101;
  assign _07707_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10100;
  assign _07708_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10011;
  assign _07709_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10010;
  assign _07710_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10001;
  assign _07711_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 5'b10000;
  assign _07712_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1111;
  assign _07713_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1110;
  assign _07714_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1101;
  assign _07715_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1100;
  assign _07716_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1011;
  assign _07717_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1010;
  assign _07718_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1001;
  assign _07719_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 4'b1000;
  assign _07720_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 3'b111;
  assign _07721_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 3'b110;
  assign _07722_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 3'b101;
  assign _07723_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 3'b100;
  assign _07724_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 2'b11;
  assign _07725_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 2'b10;
  assign _07726_ = vec_sum_050_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5566" *) 1'b1;
  function [7:0] _17195_;
    input [7:0] a;
    input [399:0] b;
    input [49:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *)
    (* parallel_case *)
    casez (s)
      50'b?????????????????????????????????????????????????1:
        _17195_ = b[7:0];
      50'b????????????????????????????????????????????????1?:
        _17195_ = b[15:8];
      50'b???????????????????????????????????????????????1??:
        _17195_ = b[23:16];
      50'b??????????????????????????????????????????????1???:
        _17195_ = b[31:24];
      50'b?????????????????????????????????????????????1????:
        _17195_ = b[39:32];
      50'b????????????????????????????????????????????1?????:
        _17195_ = b[47:40];
      50'b???????????????????????????????????????????1??????:
        _17195_ = b[55:48];
      50'b??????????????????????????????????????????1???????:
        _17195_ = b[63:56];
      50'b?????????????????????????????????????????1????????:
        _17195_ = b[71:64];
      50'b????????????????????????????????????????1?????????:
        _17195_ = b[79:72];
      50'b???????????????????????????????????????1??????????:
        _17195_ = b[87:80];
      50'b??????????????????????????????????????1???????????:
        _17195_ = b[95:88];
      50'b?????????????????????????????????????1????????????:
        _17195_ = b[103:96];
      50'b????????????????????????????????????1?????????????:
        _17195_ = b[111:104];
      50'b???????????????????????????????????1??????????????:
        _17195_ = b[119:112];
      50'b??????????????????????????????????1???????????????:
        _17195_ = b[127:120];
      50'b?????????????????????????????????1????????????????:
        _17195_ = b[135:128];
      50'b????????????????????????????????1?????????????????:
        _17195_ = b[143:136];
      50'b???????????????????????????????1??????????????????:
        _17195_ = b[151:144];
      50'b??????????????????????????????1???????????????????:
        _17195_ = b[159:152];
      50'b?????????????????????????????1????????????????????:
        _17195_ = b[167:160];
      50'b????????????????????????????1?????????????????????:
        _17195_ = b[175:168];
      50'b???????????????????????????1??????????????????????:
        _17195_ = b[183:176];
      50'b??????????????????????????1???????????????????????:
        _17195_ = b[191:184];
      50'b?????????????????????????1????????????????????????:
        _17195_ = b[199:192];
      50'b????????????????????????1?????????????????????????:
        _17195_ = b[207:200];
      50'b???????????????????????1??????????????????????????:
        _17195_ = b[215:208];
      50'b??????????????????????1???????????????????????????:
        _17195_ = b[223:216];
      50'b?????????????????????1????????????????????????????:
        _17195_ = b[231:224];
      50'b????????????????????1?????????????????????????????:
        _17195_ = b[239:232];
      50'b???????????????????1??????????????????????????????:
        _17195_ = b[247:240];
      50'b??????????????????1???????????????????????????????:
        _17195_ = b[255:248];
      50'b?????????????????1????????????????????????????????:
        _17195_ = b[263:256];
      50'b????????????????1?????????????????????????????????:
        _17195_ = b[271:264];
      50'b???????????????1??????????????????????????????????:
        _17195_ = b[279:272];
      50'b??????????????1???????????????????????????????????:
        _17195_ = b[287:280];
      50'b?????????????1????????????????????????????????????:
        _17195_ = b[295:288];
      50'b????????????1?????????????????????????????????????:
        _17195_ = b[303:296];
      50'b???????????1??????????????????????????????????????:
        _17195_ = b[311:304];
      50'b??????????1???????????????????????????????????????:
        _17195_ = b[319:312];
      50'b?????????1????????????????????????????????????????:
        _17195_ = b[327:320];
      50'b????????1?????????????????????????????????????????:
        _17195_ = b[335:328];
      50'b???????1??????????????????????????????????????????:
        _17195_ = b[343:336];
      50'b??????1???????????????????????????????????????????:
        _17195_ = b[351:344];
      50'b?????1????????????????????????????????????????????:
        _17195_ = b[359:352];
      50'b????1?????????????????????????????????????????????:
        _17195_ = b[367:360];
      50'b???1??????????????????????????????????????????????:
        _17195_ = b[375:368];
      50'b??1???????????????????????????????????????????????:
        _17195_ = b[383:376];
      50'b?1????????????????????????????????????????????????:
        _17195_ = b[391:384];
      50'b1?????????????????????????????????????????????????:
        _17195_ = b[399:392];
      default:
        _17195_ = a;
    endcase
  endfunction
  assign vec_data_049 = _17195_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384], data_d1[399:392] }, { _07776_, _07775_, _07774_, _07773_, _07772_, _07771_, _07770_, _07769_, _07768_, _07767_, _07766_, _07765_, _07764_, _07763_, _07762_, _07761_, _07760_, _07759_, _07758_, _07757_, _07756_, _07755_, _07754_, _07753_, _07752_, _07751_, _07750_, _07749_, _07748_, _07747_, _07746_, _07745_, _07744_, _07743_, _07742_, _07741_, _07740_, _07739_, _07738_, _07737_, _07736_, _07735_, _07734_, _07733_, _07732_, _07731_, _07730_, _07729_, _07728_, _07727_ });
  assign _07727_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5558|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b110010;
  assign _07728_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5557|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b110001;
  assign _07729_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5556|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b110000;
  assign _07730_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5555|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101111;
  assign _07731_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5554|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101110;
  assign _07732_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5553|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101101;
  assign _07733_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5552|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101100;
  assign _07734_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5551|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101011;
  assign _07735_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101010;
  assign _07736_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101001;
  assign _07737_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b101000;
  assign _07738_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100111;
  assign _07739_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100110;
  assign _07740_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100101;
  assign _07741_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100100;
  assign _07742_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100011;
  assign _07743_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100010;
  assign _07744_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100001;
  assign _07745_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 6'b100000;
  assign _07746_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11111;
  assign _07747_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11110;
  assign _07748_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11101;
  assign _07749_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11100;
  assign _07750_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11011;
  assign _07751_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11010;
  assign _07752_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11001;
  assign _07753_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b11000;
  assign _07754_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10111;
  assign _07755_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10110;
  assign _07756_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10101;
  assign _07757_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10100;
  assign _07758_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10011;
  assign _07759_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10010;
  assign _07760_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10001;
  assign _07761_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 5'b10000;
  assign _07762_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1111;
  assign _07763_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1110;
  assign _07764_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5521|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1101;
  assign _07765_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5520|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1100;
  assign _07766_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5519|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1011;
  assign _07767_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5518|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1010;
  assign _07768_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5517|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1001;
  assign _07769_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5516|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 4'b1000;
  assign _07770_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5515|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 3'b111;
  assign _07771_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5514|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 3'b110;
  assign _07772_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 3'b101;
  assign _07773_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 3'b100;
  assign _07774_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 2'b11;
  assign _07775_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 2'b10;
  assign _07776_ = vec_sum_049_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5508" *) 1'b1;
  function [7:0] _17246_;
    input [7:0] a;
    input [391:0] b;
    input [48:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *)
    (* parallel_case *)
    casez (s)
      49'b????????????????????????????????????????????????1:
        _17246_ = b[7:0];
      49'b???????????????????????????????????????????????1?:
        _17246_ = b[15:8];
      49'b??????????????????????????????????????????????1??:
        _17246_ = b[23:16];
      49'b?????????????????????????????????????????????1???:
        _17246_ = b[31:24];
      49'b????????????????????????????????????????????1????:
        _17246_ = b[39:32];
      49'b???????????????????????????????????????????1?????:
        _17246_ = b[47:40];
      49'b??????????????????????????????????????????1??????:
        _17246_ = b[55:48];
      49'b?????????????????????????????????????????1???????:
        _17246_ = b[63:56];
      49'b????????????????????????????????????????1????????:
        _17246_ = b[71:64];
      49'b???????????????????????????????????????1?????????:
        _17246_ = b[79:72];
      49'b??????????????????????????????????????1??????????:
        _17246_ = b[87:80];
      49'b?????????????????????????????????????1???????????:
        _17246_ = b[95:88];
      49'b????????????????????????????????????1????????????:
        _17246_ = b[103:96];
      49'b???????????????????????????????????1?????????????:
        _17246_ = b[111:104];
      49'b??????????????????????????????????1??????????????:
        _17246_ = b[119:112];
      49'b?????????????????????????????????1???????????????:
        _17246_ = b[127:120];
      49'b????????????????????????????????1????????????????:
        _17246_ = b[135:128];
      49'b???????????????????????????????1?????????????????:
        _17246_ = b[143:136];
      49'b??????????????????????????????1??????????????????:
        _17246_ = b[151:144];
      49'b?????????????????????????????1???????????????????:
        _17246_ = b[159:152];
      49'b????????????????????????????1????????????????????:
        _17246_ = b[167:160];
      49'b???????????????????????????1?????????????????????:
        _17246_ = b[175:168];
      49'b??????????????????????????1??????????????????????:
        _17246_ = b[183:176];
      49'b?????????????????????????1???????????????????????:
        _17246_ = b[191:184];
      49'b????????????????????????1????????????????????????:
        _17246_ = b[199:192];
      49'b???????????????????????1?????????????????????????:
        _17246_ = b[207:200];
      49'b??????????????????????1??????????????????????????:
        _17246_ = b[215:208];
      49'b?????????????????????1???????????????????????????:
        _17246_ = b[223:216];
      49'b????????????????????1????????????????????????????:
        _17246_ = b[231:224];
      49'b???????????????????1?????????????????????????????:
        _17246_ = b[239:232];
      49'b??????????????????1??????????????????????????????:
        _17246_ = b[247:240];
      49'b?????????????????1???????????????????????????????:
        _17246_ = b[255:248];
      49'b????????????????1????????????????????????????????:
        _17246_ = b[263:256];
      49'b???????????????1?????????????????????????????????:
        _17246_ = b[271:264];
      49'b??????????????1??????????????????????????????????:
        _17246_ = b[279:272];
      49'b?????????????1???????????????????????????????????:
        _17246_ = b[287:280];
      49'b????????????1????????????????????????????????????:
        _17246_ = b[295:288];
      49'b???????????1?????????????????????????????????????:
        _17246_ = b[303:296];
      49'b??????????1??????????????????????????????????????:
        _17246_ = b[311:304];
      49'b?????????1???????????????????????????????????????:
        _17246_ = b[319:312];
      49'b????????1????????????????????????????????????????:
        _17246_ = b[327:320];
      49'b???????1?????????????????????????????????????????:
        _17246_ = b[335:328];
      49'b??????1??????????????????????????????????????????:
        _17246_ = b[343:336];
      49'b?????1???????????????????????????????????????????:
        _17246_ = b[351:344];
      49'b????1????????????????????????????????????????????:
        _17246_ = b[359:352];
      49'b???1?????????????????????????????????????????????:
        _17246_ = b[367:360];
      49'b??1??????????????????????????????????????????????:
        _17246_ = b[375:368];
      49'b?1???????????????????????????????????????????????:
        _17246_ = b[383:376];
      49'b1????????????????????????????????????????????????:
        _17246_ = b[391:384];
      default:
        _17246_ = a;
    endcase
  endfunction
  assign vec_data_048 = _17246_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376], data_d1[391:384] }, { _07825_, _07824_, _07823_, _07822_, _07821_, _07820_, _07819_, _07818_, _07817_, _07816_, _07815_, _07814_, _07813_, _07812_, _07811_, _07810_, _07809_, _07808_, _07807_, _07806_, _07805_, _07804_, _07803_, _07802_, _07801_, _07800_, _07799_, _07798_, _07797_, _07796_, _07795_, _07794_, _07793_, _07792_, _07791_, _07790_, _07789_, _07788_, _07787_, _07786_, _07785_, _07784_, _07783_, _07782_, _07781_, _07780_, _07779_, _07778_, _07777_ });
  assign _07777_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b110001;
  assign _07778_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b110000;
  assign _07779_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101111;
  assign _07780_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101110;
  assign _07781_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101101;
  assign _07782_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101100;
  assign _07783_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101011;
  assign _07784_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101010;
  assign _07785_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101001;
  assign _07786_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b101000;
  assign _07787_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100111;
  assign _07788_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100110;
  assign _07789_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100101;
  assign _07790_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100100;
  assign _07791_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100011;
  assign _07792_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5485|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100010;
  assign _07793_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5484|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100001;
  assign _07794_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5483|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 6'b100000;
  assign _07795_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5482|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11111;
  assign _07796_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5481|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11110;
  assign _07797_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5480|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11101;
  assign _07798_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5479|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11100;
  assign _07799_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5478|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11011;
  assign _07800_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11010;
  assign _07801_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11001;
  assign _07802_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b11000;
  assign _07803_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10111;
  assign _07804_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10110;
  assign _07805_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10101;
  assign _07806_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10100;
  assign _07807_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10011;
  assign _07808_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10010;
  assign _07809_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10001;
  assign _07810_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 5'b10000;
  assign _07811_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1111;
  assign _07812_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1110;
  assign _07813_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1101;
  assign _07814_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1100;
  assign _07815_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1011;
  assign _07816_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1010;
  assign _07817_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1001;
  assign _07818_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 4'b1000;
  assign _07819_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 3'b111;
  assign _07820_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 3'b110;
  assign _07821_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 3'b101;
  assign _07822_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 3'b100;
  assign _07823_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 2'b11;
  assign _07824_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 2'b10;
  assign _07825_ = vec_sum_048_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5451" *) 1'b1;
  function [7:0] _17296_;
    input [7:0] a;
    input [383:0] b;
    input [47:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *)
    (* parallel_case *)
    casez (s)
      48'b???????????????????????????????????????????????1:
        _17296_ = b[7:0];
      48'b??????????????????????????????????????????????1?:
        _17296_ = b[15:8];
      48'b?????????????????????????????????????????????1??:
        _17296_ = b[23:16];
      48'b????????????????????????????????????????????1???:
        _17296_ = b[31:24];
      48'b???????????????????????????????????????????1????:
        _17296_ = b[39:32];
      48'b??????????????????????????????????????????1?????:
        _17296_ = b[47:40];
      48'b?????????????????????????????????????????1??????:
        _17296_ = b[55:48];
      48'b????????????????????????????????????????1???????:
        _17296_ = b[63:56];
      48'b???????????????????????????????????????1????????:
        _17296_ = b[71:64];
      48'b??????????????????????????????????????1?????????:
        _17296_ = b[79:72];
      48'b?????????????????????????????????????1??????????:
        _17296_ = b[87:80];
      48'b????????????????????????????????????1???????????:
        _17296_ = b[95:88];
      48'b???????????????????????????????????1????????????:
        _17296_ = b[103:96];
      48'b??????????????????????????????????1?????????????:
        _17296_ = b[111:104];
      48'b?????????????????????????????????1??????????????:
        _17296_ = b[119:112];
      48'b????????????????????????????????1???????????????:
        _17296_ = b[127:120];
      48'b???????????????????????????????1????????????????:
        _17296_ = b[135:128];
      48'b??????????????????????????????1?????????????????:
        _17296_ = b[143:136];
      48'b?????????????????????????????1??????????????????:
        _17296_ = b[151:144];
      48'b????????????????????????????1???????????????????:
        _17296_ = b[159:152];
      48'b???????????????????????????1????????????????????:
        _17296_ = b[167:160];
      48'b??????????????????????????1?????????????????????:
        _17296_ = b[175:168];
      48'b?????????????????????????1??????????????????????:
        _17296_ = b[183:176];
      48'b????????????????????????1???????????????????????:
        _17296_ = b[191:184];
      48'b???????????????????????1????????????????????????:
        _17296_ = b[199:192];
      48'b??????????????????????1?????????????????????????:
        _17296_ = b[207:200];
      48'b?????????????????????1??????????????????????????:
        _17296_ = b[215:208];
      48'b????????????????????1???????????????????????????:
        _17296_ = b[223:216];
      48'b???????????????????1????????????????????????????:
        _17296_ = b[231:224];
      48'b??????????????????1?????????????????????????????:
        _17296_ = b[239:232];
      48'b?????????????????1??????????????????????????????:
        _17296_ = b[247:240];
      48'b????????????????1???????????????????????????????:
        _17296_ = b[255:248];
      48'b???????????????1????????????????????????????????:
        _17296_ = b[263:256];
      48'b??????????????1?????????????????????????????????:
        _17296_ = b[271:264];
      48'b?????????????1??????????????????????????????????:
        _17296_ = b[279:272];
      48'b????????????1???????????????????????????????????:
        _17296_ = b[287:280];
      48'b???????????1????????????????????????????????????:
        _17296_ = b[295:288];
      48'b??????????1?????????????????????????????????????:
        _17296_ = b[303:296];
      48'b?????????1??????????????????????????????????????:
        _17296_ = b[311:304];
      48'b????????1???????????????????????????????????????:
        _17296_ = b[319:312];
      48'b???????1????????????????????????????????????????:
        _17296_ = b[327:320];
      48'b??????1?????????????????????????????????????????:
        _17296_ = b[335:328];
      48'b?????1??????????????????????????????????????????:
        _17296_ = b[343:336];
      48'b????1???????????????????????????????????????????:
        _17296_ = b[351:344];
      48'b???1????????????????????????????????????????????:
        _17296_ = b[359:352];
      48'b??1?????????????????????????????????????????????:
        _17296_ = b[367:360];
      48'b?1??????????????????????????????????????????????:
        _17296_ = b[375:368];
      48'b1???????????????????????????????????????????????:
        _17296_ = b[383:376];
      default:
        _17296_ = a;
    endcase
  endfunction
  assign vec_data_047 = _17296_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368], data_d1[383:376] }, { _07873_, _07872_, _07871_, _07870_, _07869_, _07868_, _07867_, _07866_, _07865_, _07864_, _07863_, _07862_, _07861_, _07860_, _07859_, _07858_, _07857_, _07856_, _07855_, _07854_, _07853_, _07852_, _07851_, _07850_, _07849_, _07848_, _07847_, _07846_, _07845_, _07844_, _07843_, _07842_, _07841_, _07840_, _07839_, _07838_, _07837_, _07836_, _07835_, _07834_, _07833_, _07832_, _07831_, _07830_, _07829_, _07828_, _07827_, _07826_ });
  assign _07826_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5443|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b110000;
  assign _07827_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101111;
  assign _07828_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101110;
  assign _07829_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101101;
  assign _07830_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101100;
  assign _07831_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101011;
  assign _07832_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101010;
  assign _07833_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101001;
  assign _07834_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b101000;
  assign _07835_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100111;
  assign _07836_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100110;
  assign _07837_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100101;
  assign _07838_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100100;
  assign _07839_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100011;
  assign _07840_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100010;
  assign _07841_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100001;
  assign _07842_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 6'b100000;
  assign _07843_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11111;
  assign _07844_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11110;
  assign _07845_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11101;
  assign _07846_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11100;
  assign _07847_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11011;
  assign _07848_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11010;
  assign _07849_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11001;
  assign _07850_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b11000;
  assign _07851_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10111;
  assign _07852_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10110;
  assign _07853_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5416|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10101;
  assign _07854_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5415|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10100;
  assign _07855_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5414|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10011;
  assign _07856_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5413|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10010;
  assign _07857_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5412|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10001;
  assign _07858_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5411|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 5'b10000;
  assign _07859_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5410|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1111;
  assign _07860_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5409|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1110;
  assign _07861_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1101;
  assign _07862_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1100;
  assign _07863_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1011;
  assign _07864_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1010;
  assign _07865_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1001;
  assign _07866_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 4'b1000;
  assign _07867_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 3'b111;
  assign _07868_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 3'b110;
  assign _07869_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 3'b101;
  assign _07870_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 3'b100;
  assign _07871_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 2'b11;
  assign _07872_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 2'b10;
  assign _07873_ = vec_sum_047_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5395" *) 1'b1;
  function [7:0] _17345_;
    input [7:0] a;
    input [375:0] b;
    input [46:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *)
    (* parallel_case *)
    casez (s)
      47'b??????????????????????????????????????????????1:
        _17345_ = b[7:0];
      47'b?????????????????????????????????????????????1?:
        _17345_ = b[15:8];
      47'b????????????????????????????????????????????1??:
        _17345_ = b[23:16];
      47'b???????????????????????????????????????????1???:
        _17345_ = b[31:24];
      47'b??????????????????????????????????????????1????:
        _17345_ = b[39:32];
      47'b?????????????????????????????????????????1?????:
        _17345_ = b[47:40];
      47'b????????????????????????????????????????1??????:
        _17345_ = b[55:48];
      47'b???????????????????????????????????????1???????:
        _17345_ = b[63:56];
      47'b??????????????????????????????????????1????????:
        _17345_ = b[71:64];
      47'b?????????????????????????????????????1?????????:
        _17345_ = b[79:72];
      47'b????????????????????????????????????1??????????:
        _17345_ = b[87:80];
      47'b???????????????????????????????????1???????????:
        _17345_ = b[95:88];
      47'b??????????????????????????????????1????????????:
        _17345_ = b[103:96];
      47'b?????????????????????????????????1?????????????:
        _17345_ = b[111:104];
      47'b????????????????????????????????1??????????????:
        _17345_ = b[119:112];
      47'b???????????????????????????????1???????????????:
        _17345_ = b[127:120];
      47'b??????????????????????????????1????????????????:
        _17345_ = b[135:128];
      47'b?????????????????????????????1?????????????????:
        _17345_ = b[143:136];
      47'b????????????????????????????1??????????????????:
        _17345_ = b[151:144];
      47'b???????????????????????????1???????????????????:
        _17345_ = b[159:152];
      47'b??????????????????????????1????????????????????:
        _17345_ = b[167:160];
      47'b?????????????????????????1?????????????????????:
        _17345_ = b[175:168];
      47'b????????????????????????1??????????????????????:
        _17345_ = b[183:176];
      47'b???????????????????????1???????????????????????:
        _17345_ = b[191:184];
      47'b??????????????????????1????????????????????????:
        _17345_ = b[199:192];
      47'b?????????????????????1?????????????????????????:
        _17345_ = b[207:200];
      47'b????????????????????1??????????????????????????:
        _17345_ = b[215:208];
      47'b???????????????????1???????????????????????????:
        _17345_ = b[223:216];
      47'b??????????????????1????????????????????????????:
        _17345_ = b[231:224];
      47'b?????????????????1?????????????????????????????:
        _17345_ = b[239:232];
      47'b????????????????1??????????????????????????????:
        _17345_ = b[247:240];
      47'b???????????????1???????????????????????????????:
        _17345_ = b[255:248];
      47'b??????????????1????????????????????????????????:
        _17345_ = b[263:256];
      47'b?????????????1?????????????????????????????????:
        _17345_ = b[271:264];
      47'b????????????1??????????????????????????????????:
        _17345_ = b[279:272];
      47'b???????????1???????????????????????????????????:
        _17345_ = b[287:280];
      47'b??????????1????????????????????????????????????:
        _17345_ = b[295:288];
      47'b?????????1?????????????????????????????????????:
        _17345_ = b[303:296];
      47'b????????1??????????????????????????????????????:
        _17345_ = b[311:304];
      47'b???????1???????????????????????????????????????:
        _17345_ = b[319:312];
      47'b??????1????????????????????????????????????????:
        _17345_ = b[327:320];
      47'b?????1?????????????????????????????????????????:
        _17345_ = b[335:328];
      47'b????1??????????????????????????????????????????:
        _17345_ = b[343:336];
      47'b???1???????????????????????????????????????????:
        _17345_ = b[351:344];
      47'b??1????????????????????????????????????????????:
        _17345_ = b[359:352];
      47'b?1?????????????????????????????????????????????:
        _17345_ = b[367:360];
      47'b1??????????????????????????????????????????????:
        _17345_ = b[375:368];
      default:
        _17345_ = a;
    endcase
  endfunction
  assign vec_data_046 = _17345_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360], data_d1[375:368] }, { _07920_, _07919_, _07918_, _07917_, _07916_, _07915_, _07914_, _07913_, _07912_, _07911_, _07910_, _07909_, _07908_, _07907_, _07906_, _07905_, _07904_, _07903_, _07902_, _07901_, _07900_, _07899_, _07898_, _07897_, _07896_, _07895_, _07894_, _07893_, _07892_, _07891_, _07890_, _07889_, _07888_, _07887_, _07886_, _07885_, _07884_, _07883_, _07882_, _07881_, _07880_, _07879_, _07878_, _07877_, _07876_, _07875_, _07874_ });
  assign _07874_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101111;
  assign _07875_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101110;
  assign _07876_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101101;
  assign _07877_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101100;
  assign _07878_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5383|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101011;
  assign _07879_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5382|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101010;
  assign _07880_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5381|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101001;
  assign _07881_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5380|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b101000;
  assign _07882_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5379|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100111;
  assign _07883_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5378|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100110;
  assign _07884_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5377|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100101;
  assign _07885_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5376|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100100;
  assign _07886_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100011;
  assign _07887_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100010;
  assign _07888_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100001;
  assign _07889_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 6'b100000;
  assign _07890_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11111;
  assign _07891_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11110;
  assign _07892_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11101;
  assign _07893_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11100;
  assign _07894_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11011;
  assign _07895_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11010;
  assign _07896_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11001;
  assign _07897_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b11000;
  assign _07898_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10111;
  assign _07899_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10110;
  assign _07900_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10101;
  assign _07901_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10100;
  assign _07902_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10011;
  assign _07903_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10010;
  assign _07904_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10001;
  assign _07905_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 5'b10000;
  assign _07906_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1111;
  assign _07907_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1110;
  assign _07908_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1101;
  assign _07909_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1100;
  assign _07910_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5351|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1011;
  assign _07911_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5350|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1010;
  assign _07912_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5349|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1001;
  assign _07913_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5348|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 4'b1000;
  assign _07914_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5347|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 3'b111;
  assign _07915_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5346|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 3'b110;
  assign _07916_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5345|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 3'b101;
  assign _07917_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5344|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 3'b100;
  assign _07918_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 2'b11;
  assign _07919_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 2'b10;
  assign _07920_ = vec_sum_046_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5340" *) 1'b1;
  function [7:0] _17393_;
    input [7:0] a;
    input [367:0] b;
    input [45:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *)
    (* parallel_case *)
    casez (s)
      46'b?????????????????????????????????????????????1:
        _17393_ = b[7:0];
      46'b????????????????????????????????????????????1?:
        _17393_ = b[15:8];
      46'b???????????????????????????????????????????1??:
        _17393_ = b[23:16];
      46'b??????????????????????????????????????????1???:
        _17393_ = b[31:24];
      46'b?????????????????????????????????????????1????:
        _17393_ = b[39:32];
      46'b????????????????????????????????????????1?????:
        _17393_ = b[47:40];
      46'b???????????????????????????????????????1??????:
        _17393_ = b[55:48];
      46'b??????????????????????????????????????1???????:
        _17393_ = b[63:56];
      46'b?????????????????????????????????????1????????:
        _17393_ = b[71:64];
      46'b????????????????????????????????????1?????????:
        _17393_ = b[79:72];
      46'b???????????????????????????????????1??????????:
        _17393_ = b[87:80];
      46'b??????????????????????????????????1???????????:
        _17393_ = b[95:88];
      46'b?????????????????????????????????1????????????:
        _17393_ = b[103:96];
      46'b????????????????????????????????1?????????????:
        _17393_ = b[111:104];
      46'b???????????????????????????????1??????????????:
        _17393_ = b[119:112];
      46'b??????????????????????????????1???????????????:
        _17393_ = b[127:120];
      46'b?????????????????????????????1????????????????:
        _17393_ = b[135:128];
      46'b????????????????????????????1?????????????????:
        _17393_ = b[143:136];
      46'b???????????????????????????1??????????????????:
        _17393_ = b[151:144];
      46'b??????????????????????????1???????????????????:
        _17393_ = b[159:152];
      46'b?????????????????????????1????????????????????:
        _17393_ = b[167:160];
      46'b????????????????????????1?????????????????????:
        _17393_ = b[175:168];
      46'b???????????????????????1??????????????????????:
        _17393_ = b[183:176];
      46'b??????????????????????1???????????????????????:
        _17393_ = b[191:184];
      46'b?????????????????????1????????????????????????:
        _17393_ = b[199:192];
      46'b????????????????????1?????????????????????????:
        _17393_ = b[207:200];
      46'b???????????????????1??????????????????????????:
        _17393_ = b[215:208];
      46'b??????????????????1???????????????????????????:
        _17393_ = b[223:216];
      46'b?????????????????1????????????????????????????:
        _17393_ = b[231:224];
      46'b????????????????1?????????????????????????????:
        _17393_ = b[239:232];
      46'b???????????????1??????????????????????????????:
        _17393_ = b[247:240];
      46'b??????????????1???????????????????????????????:
        _17393_ = b[255:248];
      46'b?????????????1????????????????????????????????:
        _17393_ = b[263:256];
      46'b????????????1?????????????????????????????????:
        _17393_ = b[271:264];
      46'b???????????1??????????????????????????????????:
        _17393_ = b[279:272];
      46'b??????????1???????????????????????????????????:
        _17393_ = b[287:280];
      46'b?????????1????????????????????????????????????:
        _17393_ = b[295:288];
      46'b????????1?????????????????????????????????????:
        _17393_ = b[303:296];
      46'b???????1??????????????????????????????????????:
        _17393_ = b[311:304];
      46'b??????1???????????????????????????????????????:
        _17393_ = b[319:312];
      46'b?????1????????????????????????????????????????:
        _17393_ = b[327:320];
      46'b????1?????????????????????????????????????????:
        _17393_ = b[335:328];
      46'b???1??????????????????????????????????????????:
        _17393_ = b[343:336];
      46'b??1???????????????????????????????????????????:
        _17393_ = b[351:344];
      46'b?1????????????????????????????????????????????:
        _17393_ = b[359:352];
      46'b1?????????????????????????????????????????????:
        _17393_ = b[367:360];
      default:
        _17393_ = a;
    endcase
  endfunction
  assign vec_data_045 = _17393_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352], data_d1[367:360] }, { _07966_, _07965_, _07964_, _07963_, _07962_, _07961_, _07960_, _07959_, _07958_, _07957_, _07956_, _07955_, _07954_, _07953_, _07952_, _07951_, _07950_, _07949_, _07948_, _07947_, _07946_, _07945_, _07944_, _07943_, _07942_, _07941_, _07940_, _07939_, _07938_, _07937_, _07936_, _07935_, _07934_, _07933_, _07932_, _07931_, _07930_, _07929_, _07928_, _07927_, _07926_, _07925_, _07924_, _07923_, _07922_, _07921_ });
  assign _07921_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101110;
  assign _07922_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101101;
  assign _07923_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101100;
  assign _07924_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101011;
  assign _07925_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101010;
  assign _07926_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101001;
  assign _07927_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b101000;
  assign _07928_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100111;
  assign _07929_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100110;
  assign _07930_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100101;
  assign _07931_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100100;
  assign _07932_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100011;
  assign _07933_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5320|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100010;
  assign _07934_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5319|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100001;
  assign _07935_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5318|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 6'b100000;
  assign _07936_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5317|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11111;
  assign _07937_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5316|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11110;
  assign _07938_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5315|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11101;
  assign _07939_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5314|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11100;
  assign _07940_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5313|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11011;
  assign _07941_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11010;
  assign _07942_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11001;
  assign _07943_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b11000;
  assign _07944_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10111;
  assign _07945_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10110;
  assign _07946_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10101;
  assign _07947_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10100;
  assign _07948_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10011;
  assign _07949_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10010;
  assign _07950_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10001;
  assign _07951_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 5'b10000;
  assign _07952_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1111;
  assign _07953_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1110;
  assign _07954_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1101;
  assign _07955_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1100;
  assign _07956_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1011;
  assign _07957_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1010;
  assign _07958_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1001;
  assign _07959_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 4'b1000;
  assign _07960_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 3'b111;
  assign _07961_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 3'b110;
  assign _07962_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 3'b101;
  assign _07963_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5290|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 3'b100;
  assign _07964_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5289|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 2'b11;
  assign _07965_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5288|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 2'b10;
  assign _07966_ = vec_sum_045_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5287|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5286" *) 1'b1;
  function [7:0] _17440_;
    input [7:0] a;
    input [359:0] b;
    input [44:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *)
    (* parallel_case *)
    casez (s)
      45'b????????????????????????????????????????????1:
        _17440_ = b[7:0];
      45'b???????????????????????????????????????????1?:
        _17440_ = b[15:8];
      45'b??????????????????????????????????????????1??:
        _17440_ = b[23:16];
      45'b?????????????????????????????????????????1???:
        _17440_ = b[31:24];
      45'b????????????????????????????????????????1????:
        _17440_ = b[39:32];
      45'b???????????????????????????????????????1?????:
        _17440_ = b[47:40];
      45'b??????????????????????????????????????1??????:
        _17440_ = b[55:48];
      45'b?????????????????????????????????????1???????:
        _17440_ = b[63:56];
      45'b????????????????????????????????????1????????:
        _17440_ = b[71:64];
      45'b???????????????????????????????????1?????????:
        _17440_ = b[79:72];
      45'b??????????????????????????????????1??????????:
        _17440_ = b[87:80];
      45'b?????????????????????????????????1???????????:
        _17440_ = b[95:88];
      45'b????????????????????????????????1????????????:
        _17440_ = b[103:96];
      45'b???????????????????????????????1?????????????:
        _17440_ = b[111:104];
      45'b??????????????????????????????1??????????????:
        _17440_ = b[119:112];
      45'b?????????????????????????????1???????????????:
        _17440_ = b[127:120];
      45'b????????????????????????????1????????????????:
        _17440_ = b[135:128];
      45'b???????????????????????????1?????????????????:
        _17440_ = b[143:136];
      45'b??????????????????????????1??????????????????:
        _17440_ = b[151:144];
      45'b?????????????????????????1???????????????????:
        _17440_ = b[159:152];
      45'b????????????????????????1????????????????????:
        _17440_ = b[167:160];
      45'b???????????????????????1?????????????????????:
        _17440_ = b[175:168];
      45'b??????????????????????1??????????????????????:
        _17440_ = b[183:176];
      45'b?????????????????????1???????????????????????:
        _17440_ = b[191:184];
      45'b????????????????????1????????????????????????:
        _17440_ = b[199:192];
      45'b???????????????????1?????????????????????????:
        _17440_ = b[207:200];
      45'b??????????????????1??????????????????????????:
        _17440_ = b[215:208];
      45'b?????????????????1???????????????????????????:
        _17440_ = b[223:216];
      45'b????????????????1????????????????????????????:
        _17440_ = b[231:224];
      45'b???????????????1?????????????????????????????:
        _17440_ = b[239:232];
      45'b??????????????1??????????????????????????????:
        _17440_ = b[247:240];
      45'b?????????????1???????????????????????????????:
        _17440_ = b[255:248];
      45'b????????????1????????????????????????????????:
        _17440_ = b[263:256];
      45'b???????????1?????????????????????????????????:
        _17440_ = b[271:264];
      45'b??????????1??????????????????????????????????:
        _17440_ = b[279:272];
      45'b?????????1???????????????????????????????????:
        _17440_ = b[287:280];
      45'b????????1????????????????????????????????????:
        _17440_ = b[295:288];
      45'b???????1?????????????????????????????????????:
        _17440_ = b[303:296];
      45'b??????1??????????????????????????????????????:
        _17440_ = b[311:304];
      45'b?????1???????????????????????????????????????:
        _17440_ = b[319:312];
      45'b????1????????????????????????????????????????:
        _17440_ = b[327:320];
      45'b???1?????????????????????????????????????????:
        _17440_ = b[335:328];
      45'b??1??????????????????????????????????????????:
        _17440_ = b[343:336];
      45'b?1???????????????????????????????????????????:
        _17440_ = b[351:344];
      45'b1????????????????????????????????????????????:
        _17440_ = b[359:352];
      default:
        _17440_ = a;
    endcase
  endfunction
  assign vec_data_044 = _17440_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344], data_d1[359:352] }, { _08011_, _08010_, _08009_, _08008_, _08007_, _08006_, _08005_, _08004_, _08003_, _08002_, _08001_, _08000_, _07999_, _07998_, _07997_, _07996_, _07995_, _07994_, _07993_, _07992_, _07991_, _07990_, _07989_, _07988_, _07987_, _07986_, _07985_, _07984_, _07983_, _07982_, _07981_, _07980_, _07979_, _07978_, _07977_, _07976_, _07975_, _07974_, _07973_, _07972_, _07971_, _07970_, _07969_, _07968_, _07967_ });
  assign _07967_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101101;
  assign _07968_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101100;
  assign _07969_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101011;
  assign _07970_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101010;
  assign _07971_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101001;
  assign _07972_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b101000;
  assign _07973_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100111;
  assign _07974_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100110;
  assign _07975_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100101;
  assign _07976_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100100;
  assign _07977_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100011;
  assign _07978_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100010;
  assign _07979_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100001;
  assign _07980_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 6'b100000;
  assign _07981_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11111;
  assign _07982_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11110;
  assign _07983_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11101;
  assign _07984_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5261|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11100;
  assign _07985_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5260|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11011;
  assign _07986_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5259|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11010;
  assign _07987_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5258|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11001;
  assign _07988_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5257|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b11000;
  assign _07989_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5256|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10111;
  assign _07990_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5255|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10110;
  assign _07991_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5254|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10101;
  assign _07992_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10100;
  assign _07993_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10011;
  assign _07994_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10010;
  assign _07995_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10001;
  assign _07996_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 5'b10000;
  assign _07997_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1111;
  assign _07998_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1110;
  assign _07999_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1101;
  assign _08000_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1100;
  assign _08001_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1011;
  assign _08002_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1010;
  assign _08003_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1001;
  assign _08004_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 4'b1000;
  assign _08005_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 3'b111;
  assign _08006_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 3'b110;
  assign _08007_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 3'b101;
  assign _08008_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 3'b100;
  assign _08009_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 2'b11;
  assign _08010_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 2'b10;
  assign _08011_ = vec_sum_044_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5233" *) 1'b1;
  function [7:0] _17486_;
    input [7:0] a;
    input [351:0] b;
    input [43:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *)
    (* parallel_case *)
    casez (s)
      44'b???????????????????????????????????????????1:
        _17486_ = b[7:0];
      44'b??????????????????????????????????????????1?:
        _17486_ = b[15:8];
      44'b?????????????????????????????????????????1??:
        _17486_ = b[23:16];
      44'b????????????????????????????????????????1???:
        _17486_ = b[31:24];
      44'b???????????????????????????????????????1????:
        _17486_ = b[39:32];
      44'b??????????????????????????????????????1?????:
        _17486_ = b[47:40];
      44'b?????????????????????????????????????1??????:
        _17486_ = b[55:48];
      44'b????????????????????????????????????1???????:
        _17486_ = b[63:56];
      44'b???????????????????????????????????1????????:
        _17486_ = b[71:64];
      44'b??????????????????????????????????1?????????:
        _17486_ = b[79:72];
      44'b?????????????????????????????????1??????????:
        _17486_ = b[87:80];
      44'b????????????????????????????????1???????????:
        _17486_ = b[95:88];
      44'b???????????????????????????????1????????????:
        _17486_ = b[103:96];
      44'b??????????????????????????????1?????????????:
        _17486_ = b[111:104];
      44'b?????????????????????????????1??????????????:
        _17486_ = b[119:112];
      44'b????????????????????????????1???????????????:
        _17486_ = b[127:120];
      44'b???????????????????????????1????????????????:
        _17486_ = b[135:128];
      44'b??????????????????????????1?????????????????:
        _17486_ = b[143:136];
      44'b?????????????????????????1??????????????????:
        _17486_ = b[151:144];
      44'b????????????????????????1???????????????????:
        _17486_ = b[159:152];
      44'b???????????????????????1????????????????????:
        _17486_ = b[167:160];
      44'b??????????????????????1?????????????????????:
        _17486_ = b[175:168];
      44'b?????????????????????1??????????????????????:
        _17486_ = b[183:176];
      44'b????????????????????1???????????????????????:
        _17486_ = b[191:184];
      44'b???????????????????1????????????????????????:
        _17486_ = b[199:192];
      44'b??????????????????1?????????????????????????:
        _17486_ = b[207:200];
      44'b?????????????????1??????????????????????????:
        _17486_ = b[215:208];
      44'b????????????????1???????????????????????????:
        _17486_ = b[223:216];
      44'b???????????????1????????????????????????????:
        _17486_ = b[231:224];
      44'b??????????????1?????????????????????????????:
        _17486_ = b[239:232];
      44'b?????????????1??????????????????????????????:
        _17486_ = b[247:240];
      44'b????????????1???????????????????????????????:
        _17486_ = b[255:248];
      44'b???????????1????????????????????????????????:
        _17486_ = b[263:256];
      44'b??????????1?????????????????????????????????:
        _17486_ = b[271:264];
      44'b?????????1??????????????????????????????????:
        _17486_ = b[279:272];
      44'b????????1???????????????????????????????????:
        _17486_ = b[287:280];
      44'b???????1????????????????????????????????????:
        _17486_ = b[295:288];
      44'b??????1?????????????????????????????????????:
        _17486_ = b[303:296];
      44'b?????1??????????????????????????????????????:
        _17486_ = b[311:304];
      44'b????1???????????????????????????????????????:
        _17486_ = b[319:312];
      44'b???1????????????????????????????????????????:
        _17486_ = b[327:320];
      44'b??1?????????????????????????????????????????:
        _17486_ = b[335:328];
      44'b?1??????????????????????????????????????????:
        _17486_ = b[343:336];
      44'b1???????????????????????????????????????????:
        _17486_ = b[351:344];
      default:
        _17486_ = a;
    endcase
  endfunction
  assign vec_data_043 = _17486_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336], data_d1[351:344] }, { _08055_, _08054_, _08053_, _08052_, _08051_, _08050_, _08049_, _08048_, _08047_, _08046_, _08045_, _08044_, _08043_, _08042_, _08041_, _08040_, _08039_, _08038_, _08037_, _08036_, _08035_, _08034_, _08033_, _08032_, _08031_, _08030_, _08029_, _08028_, _08027_, _08026_, _08025_, _08024_, _08023_, _08022_, _08021_, _08020_, _08019_, _08018_, _08017_, _08016_, _08015_, _08014_, _08013_, _08012_ });
  assign _08012_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b101100;
  assign _08013_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b101011;
  assign _08014_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b101010;
  assign _08015_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b101001;
  assign _08016_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b101000;
  assign _08017_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100111;
  assign _08018_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100110;
  assign _08019_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100101;
  assign _08020_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100100;
  assign _08021_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100011;
  assign _08022_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100010;
  assign _08023_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100001;
  assign _08024_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 6'b100000;
  assign _08025_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11111;
  assign _08026_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11110;
  assign _08027_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11101;
  assign _08028_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11100;
  assign _08029_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11011;
  assign _08030_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11010;
  assign _08031_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5206|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11001;
  assign _08032_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5205|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b11000;
  assign _08033_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5204|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10111;
  assign _08034_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5203|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10110;
  assign _08035_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5202|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10101;
  assign _08036_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5201|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10100;
  assign _08037_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5200|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10011;
  assign _08038_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5199|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10010;
  assign _08039_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10001;
  assign _08040_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 5'b10000;
  assign _08041_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1111;
  assign _08042_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1110;
  assign _08043_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1101;
  assign _08044_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1100;
  assign _08045_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1011;
  assign _08046_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1010;
  assign _08047_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1001;
  assign _08048_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 4'b1000;
  assign _08049_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 3'b111;
  assign _08050_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 3'b110;
  assign _08051_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 3'b101;
  assign _08052_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 3'b100;
  assign _08053_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 2'b11;
  assign _08054_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 2'b10;
  assign _08055_ = vec_sum_043_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5181" *) 1'b1;
  function [7:0] _17531_;
    input [7:0] a;
    input [343:0] b;
    input [42:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *)
    (* parallel_case *)
    casez (s)
      43'b??????????????????????????????????????????1:
        _17531_ = b[7:0];
      43'b?????????????????????????????????????????1?:
        _17531_ = b[15:8];
      43'b????????????????????????????????????????1??:
        _17531_ = b[23:16];
      43'b???????????????????????????????????????1???:
        _17531_ = b[31:24];
      43'b??????????????????????????????????????1????:
        _17531_ = b[39:32];
      43'b?????????????????????????????????????1?????:
        _17531_ = b[47:40];
      43'b????????????????????????????????????1??????:
        _17531_ = b[55:48];
      43'b???????????????????????????????????1???????:
        _17531_ = b[63:56];
      43'b??????????????????????????????????1????????:
        _17531_ = b[71:64];
      43'b?????????????????????????????????1?????????:
        _17531_ = b[79:72];
      43'b????????????????????????????????1??????????:
        _17531_ = b[87:80];
      43'b???????????????????????????????1???????????:
        _17531_ = b[95:88];
      43'b??????????????????????????????1????????????:
        _17531_ = b[103:96];
      43'b?????????????????????????????1?????????????:
        _17531_ = b[111:104];
      43'b????????????????????????????1??????????????:
        _17531_ = b[119:112];
      43'b???????????????????????????1???????????????:
        _17531_ = b[127:120];
      43'b??????????????????????????1????????????????:
        _17531_ = b[135:128];
      43'b?????????????????????????1?????????????????:
        _17531_ = b[143:136];
      43'b????????????????????????1??????????????????:
        _17531_ = b[151:144];
      43'b???????????????????????1???????????????????:
        _17531_ = b[159:152];
      43'b??????????????????????1????????????????????:
        _17531_ = b[167:160];
      43'b?????????????????????1?????????????????????:
        _17531_ = b[175:168];
      43'b????????????????????1??????????????????????:
        _17531_ = b[183:176];
      43'b???????????????????1???????????????????????:
        _17531_ = b[191:184];
      43'b??????????????????1????????????????????????:
        _17531_ = b[199:192];
      43'b?????????????????1?????????????????????????:
        _17531_ = b[207:200];
      43'b????????????????1??????????????????????????:
        _17531_ = b[215:208];
      43'b???????????????1???????????????????????????:
        _17531_ = b[223:216];
      43'b??????????????1????????????????????????????:
        _17531_ = b[231:224];
      43'b?????????????1?????????????????????????????:
        _17531_ = b[239:232];
      43'b????????????1??????????????????????????????:
        _17531_ = b[247:240];
      43'b???????????1???????????????????????????????:
        _17531_ = b[255:248];
      43'b??????????1????????????????????????????????:
        _17531_ = b[263:256];
      43'b?????????1?????????????????????????????????:
        _17531_ = b[271:264];
      43'b????????1??????????????????????????????????:
        _17531_ = b[279:272];
      43'b???????1???????????????????????????????????:
        _17531_ = b[287:280];
      43'b??????1????????????????????????????????????:
        _17531_ = b[295:288];
      43'b?????1?????????????????????????????????????:
        _17531_ = b[303:296];
      43'b????1??????????????????????????????????????:
        _17531_ = b[311:304];
      43'b???1???????????????????????????????????????:
        _17531_ = b[319:312];
      43'b??1????????????????????????????????????????:
        _17531_ = b[327:320];
      43'b?1?????????????????????????????????????????:
        _17531_ = b[335:328];
      43'b1??????????????????????????????????????????:
        _17531_ = b[343:336];
      default:
        _17531_ = a;
    endcase
  endfunction
  assign vec_data_042 = _17531_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328], data_d1[343:336] }, { _08098_, _08097_, _08096_, _08095_, _08094_, _08093_, _08092_, _08091_, _08090_, _08089_, _08088_, _08087_, _08086_, _08085_, _08084_, _08083_, _08082_, _08081_, _08080_, _08079_, _08078_, _08077_, _08076_, _08075_, _08074_, _08073_, _08072_, _08071_, _08070_, _08069_, _08068_, _08067_, _08066_, _08065_, _08064_, _08063_, _08062_, _08061_, _08060_, _08059_, _08058_, _08057_, _08056_ });
  assign _08056_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5173|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b101011;
  assign _08057_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b101010;
  assign _08058_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b101001;
  assign _08059_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b101000;
  assign _08060_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100111;
  assign _08061_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100110;
  assign _08062_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100101;
  assign _08063_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100100;
  assign _08064_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100011;
  assign _08065_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100010;
  assign _08066_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100001;
  assign _08067_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 6'b100000;
  assign _08068_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11111;
  assign _08069_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11110;
  assign _08070_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11101;
  assign _08071_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11100;
  assign _08072_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11011;
  assign _08073_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11010;
  assign _08074_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5155|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11001;
  assign _08075_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5154|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b11000;
  assign _08076_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5153|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10111;
  assign _08077_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5152|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10110;
  assign _08078_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5151|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10101;
  assign _08079_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5150|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10100;
  assign _08080_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5149|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10011;
  assign _08081_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5148|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10010;
  assign _08082_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10001;
  assign _08083_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 5'b10000;
  assign _08084_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1111;
  assign _08085_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1110;
  assign _08086_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1101;
  assign _08087_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1100;
  assign _08088_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1011;
  assign _08089_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1010;
  assign _08090_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1001;
  assign _08091_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 4'b1000;
  assign _08092_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 3'b111;
  assign _08093_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 3'b110;
  assign _08094_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 3'b101;
  assign _08095_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 3'b100;
  assign _08096_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 2'b11;
  assign _08097_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 2'b10;
  assign _08098_ = vec_sum_042_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5131|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5130" *) 1'b1;
  function [7:0] _17575_;
    input [7:0] a;
    input [335:0] b;
    input [41:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *)
    (* parallel_case *)
    casez (s)
      42'b?????????????????????????????????????????1:
        _17575_ = b[7:0];
      42'b????????????????????????????????????????1?:
        _17575_ = b[15:8];
      42'b???????????????????????????????????????1??:
        _17575_ = b[23:16];
      42'b??????????????????????????????????????1???:
        _17575_ = b[31:24];
      42'b?????????????????????????????????????1????:
        _17575_ = b[39:32];
      42'b????????????????????????????????????1?????:
        _17575_ = b[47:40];
      42'b???????????????????????????????????1??????:
        _17575_ = b[55:48];
      42'b??????????????????????????????????1???????:
        _17575_ = b[63:56];
      42'b?????????????????????????????????1????????:
        _17575_ = b[71:64];
      42'b????????????????????????????????1?????????:
        _17575_ = b[79:72];
      42'b???????????????????????????????1??????????:
        _17575_ = b[87:80];
      42'b??????????????????????????????1???????????:
        _17575_ = b[95:88];
      42'b?????????????????????????????1????????????:
        _17575_ = b[103:96];
      42'b????????????????????????????1?????????????:
        _17575_ = b[111:104];
      42'b???????????????????????????1??????????????:
        _17575_ = b[119:112];
      42'b??????????????????????????1???????????????:
        _17575_ = b[127:120];
      42'b?????????????????????????1????????????????:
        _17575_ = b[135:128];
      42'b????????????????????????1?????????????????:
        _17575_ = b[143:136];
      42'b???????????????????????1??????????????????:
        _17575_ = b[151:144];
      42'b??????????????????????1???????????????????:
        _17575_ = b[159:152];
      42'b?????????????????????1????????????????????:
        _17575_ = b[167:160];
      42'b????????????????????1?????????????????????:
        _17575_ = b[175:168];
      42'b???????????????????1??????????????????????:
        _17575_ = b[183:176];
      42'b??????????????????1???????????????????????:
        _17575_ = b[191:184];
      42'b?????????????????1????????????????????????:
        _17575_ = b[199:192];
      42'b????????????????1?????????????????????????:
        _17575_ = b[207:200];
      42'b???????????????1??????????????????????????:
        _17575_ = b[215:208];
      42'b??????????????1???????????????????????????:
        _17575_ = b[223:216];
      42'b?????????????1????????????????????????????:
        _17575_ = b[231:224];
      42'b????????????1?????????????????????????????:
        _17575_ = b[239:232];
      42'b???????????1??????????????????????????????:
        _17575_ = b[247:240];
      42'b??????????1???????????????????????????????:
        _17575_ = b[255:248];
      42'b?????????1????????????????????????????????:
        _17575_ = b[263:256];
      42'b????????1?????????????????????????????????:
        _17575_ = b[271:264];
      42'b???????1??????????????????????????????????:
        _17575_ = b[279:272];
      42'b??????1???????????????????????????????????:
        _17575_ = b[287:280];
      42'b?????1????????????????????????????????????:
        _17575_ = b[295:288];
      42'b????1?????????????????????????????????????:
        _17575_ = b[303:296];
      42'b???1??????????????????????????????????????:
        _17575_ = b[311:304];
      42'b??1???????????????????????????????????????:
        _17575_ = b[319:312];
      42'b?1????????????????????????????????????????:
        _17575_ = b[327:320];
      42'b1?????????????????????????????????????????:
        _17575_ = b[335:328];
      default:
        _17575_ = a;
    endcase
  endfunction
  assign vec_data_041 = _17575_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320], data_d1[335:328] }, { _08140_, _08139_, _08138_, _08137_, _08136_, _08135_, _08134_, _08133_, _08132_, _08131_, _08130_, _08129_, _08128_, _08127_, _08126_, _08125_, _08124_, _08123_, _08122_, _08121_, _08120_, _08119_, _08118_, _08117_, _08116_, _08115_, _08114_, _08113_, _08112_, _08111_, _08110_, _08109_, _08108_, _08107_, _08106_, _08105_, _08104_, _08103_, _08102_, _08101_, _08100_, _08099_ });
  assign _08099_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b101010;
  assign _08100_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b101001;
  assign _08101_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b101000;
  assign _08102_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100111;
  assign _08103_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100110;
  assign _08104_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100101;
  assign _08105_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100100;
  assign _08106_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100011;
  assign _08107_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100010;
  assign _08108_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100001;
  assign _08109_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 6'b100000;
  assign _08110_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11111;
  assign _08111_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11110;
  assign _08112_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11101;
  assign _08113_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5108|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11100;
  assign _08114_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5107|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11011;
  assign _08115_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5106|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11010;
  assign _08116_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5105|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11001;
  assign _08117_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5104|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b11000;
  assign _08118_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5103|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10111;
  assign _08119_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5102|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10110;
  assign _08120_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5101|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10101;
  assign _08121_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10100;
  assign _08122_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10011;
  assign _08123_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10010;
  assign _08124_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10001;
  assign _08125_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 5'b10000;
  assign _08126_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1111;
  assign _08127_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1110;
  assign _08128_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1101;
  assign _08129_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1100;
  assign _08130_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1011;
  assign _08131_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1010;
  assign _08132_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1001;
  assign _08133_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 4'b1000;
  assign _08134_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 3'b111;
  assign _08135_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5086|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 3'b110;
  assign _08136_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5085|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 3'b101;
  assign _08137_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5084|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 3'b100;
  assign _08138_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5083|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 2'b11;
  assign _08139_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5082|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 2'b10;
  assign _08140_ = vec_sum_041_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5081|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5080" *) 1'b1;
  function [7:0] _17618_;
    input [7:0] a;
    input [327:0] b;
    input [40:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *)
    (* parallel_case *)
    casez (s)
      41'b????????????????????????????????????????1:
        _17618_ = b[7:0];
      41'b???????????????????????????????????????1?:
        _17618_ = b[15:8];
      41'b??????????????????????????????????????1??:
        _17618_ = b[23:16];
      41'b?????????????????????????????????????1???:
        _17618_ = b[31:24];
      41'b????????????????????????????????????1????:
        _17618_ = b[39:32];
      41'b???????????????????????????????????1?????:
        _17618_ = b[47:40];
      41'b??????????????????????????????????1??????:
        _17618_ = b[55:48];
      41'b?????????????????????????????????1???????:
        _17618_ = b[63:56];
      41'b????????????????????????????????1????????:
        _17618_ = b[71:64];
      41'b???????????????????????????????1?????????:
        _17618_ = b[79:72];
      41'b??????????????????????????????1??????????:
        _17618_ = b[87:80];
      41'b?????????????????????????????1???????????:
        _17618_ = b[95:88];
      41'b????????????????????????????1????????????:
        _17618_ = b[103:96];
      41'b???????????????????????????1?????????????:
        _17618_ = b[111:104];
      41'b??????????????????????????1??????????????:
        _17618_ = b[119:112];
      41'b?????????????????????????1???????????????:
        _17618_ = b[127:120];
      41'b????????????????????????1????????????????:
        _17618_ = b[135:128];
      41'b???????????????????????1?????????????????:
        _17618_ = b[143:136];
      41'b??????????????????????1??????????????????:
        _17618_ = b[151:144];
      41'b?????????????????????1???????????????????:
        _17618_ = b[159:152];
      41'b????????????????????1????????????????????:
        _17618_ = b[167:160];
      41'b???????????????????1?????????????????????:
        _17618_ = b[175:168];
      41'b??????????????????1??????????????????????:
        _17618_ = b[183:176];
      41'b?????????????????1???????????????????????:
        _17618_ = b[191:184];
      41'b????????????????1????????????????????????:
        _17618_ = b[199:192];
      41'b???????????????1?????????????????????????:
        _17618_ = b[207:200];
      41'b??????????????1??????????????????????????:
        _17618_ = b[215:208];
      41'b?????????????1???????????????????????????:
        _17618_ = b[223:216];
      41'b????????????1????????????????????????????:
        _17618_ = b[231:224];
      41'b???????????1?????????????????????????????:
        _17618_ = b[239:232];
      41'b??????????1??????????????????????????????:
        _17618_ = b[247:240];
      41'b?????????1???????????????????????????????:
        _17618_ = b[255:248];
      41'b????????1????????????????????????????????:
        _17618_ = b[263:256];
      41'b???????1?????????????????????????????????:
        _17618_ = b[271:264];
      41'b??????1??????????????????????????????????:
        _17618_ = b[279:272];
      41'b?????1???????????????????????????????????:
        _17618_ = b[287:280];
      41'b????1????????????????????????????????????:
        _17618_ = b[295:288];
      41'b???1?????????????????????????????????????:
        _17618_ = b[303:296];
      41'b??1??????????????????????????????????????:
        _17618_ = b[311:304];
      41'b?1???????????????????????????????????????:
        _17618_ = b[319:312];
      41'b1????????????????????????????????????????:
        _17618_ = b[327:320];
      default:
        _17618_ = a;
    endcase
  endfunction
  assign vec_data_040 = _17618_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312], data_d1[327:320] }, { _08181_, _08180_, _08179_, _08178_, _08177_, _08176_, _08175_, _08174_, _08173_, _08172_, _08171_, _08170_, _08169_, _08168_, _08167_, _08166_, _08165_, _08164_, _08163_, _08162_, _08161_, _08160_, _08159_, _08158_, _08157_, _08156_, _08155_, _08154_, _08153_, _08152_, _08151_, _08150_, _08149_, _08148_, _08147_, _08146_, _08145_, _08144_, _08143_, _08142_, _08141_ });
  assign _08141_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b101001;
  assign _08142_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b101000;
  assign _08143_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100111;
  assign _08144_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100110;
  assign _08145_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100101;
  assign _08146_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100100;
  assign _08147_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100011;
  assign _08148_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5065|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100010;
  assign _08149_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5064|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100001;
  assign _08150_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5063|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 6'b100000;
  assign _08151_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5062|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11111;
  assign _08152_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5061|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11110;
  assign _08153_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5060|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11101;
  assign _08154_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5059|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11100;
  assign _08155_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5058|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11011;
  assign _08156_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11010;
  assign _08157_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11001;
  assign _08158_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b11000;
  assign _08159_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10111;
  assign _08160_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10110;
  assign _08161_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10101;
  assign _08162_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10100;
  assign _08163_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10011;
  assign _08164_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10010;
  assign _08165_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10001;
  assign _08166_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 5'b10000;
  assign _08167_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1111;
  assign _08168_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5045|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1110;
  assign _08169_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5044|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1101;
  assign _08170_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5043|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1100;
  assign _08171_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5042|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1011;
  assign _08172_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5041|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1010;
  assign _08173_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5040|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1001;
  assign _08174_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5039|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 4'b1000;
  assign _08175_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5038|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 3'b111;
  assign _08176_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 3'b110;
  assign _08177_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 3'b101;
  assign _08178_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 3'b100;
  assign _08179_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 2'b11;
  assign _08180_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 2'b10;
  assign _08181_ = vec_sum_040_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5031" *) 1'b1;
  function [7:0] _17660_;
    input [7:0] a;
    input [319:0] b;
    input [39:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *)
    (* parallel_case *)
    casez (s)
      40'b???????????????????????????????????????1:
        _17660_ = b[7:0];
      40'b??????????????????????????????????????1?:
        _17660_ = b[15:8];
      40'b?????????????????????????????????????1??:
        _17660_ = b[23:16];
      40'b????????????????????????????????????1???:
        _17660_ = b[31:24];
      40'b???????????????????????????????????1????:
        _17660_ = b[39:32];
      40'b??????????????????????????????????1?????:
        _17660_ = b[47:40];
      40'b?????????????????????????????????1??????:
        _17660_ = b[55:48];
      40'b????????????????????????????????1???????:
        _17660_ = b[63:56];
      40'b???????????????????????????????1????????:
        _17660_ = b[71:64];
      40'b??????????????????????????????1?????????:
        _17660_ = b[79:72];
      40'b?????????????????????????????1??????????:
        _17660_ = b[87:80];
      40'b????????????????????????????1???????????:
        _17660_ = b[95:88];
      40'b???????????????????????????1????????????:
        _17660_ = b[103:96];
      40'b??????????????????????????1?????????????:
        _17660_ = b[111:104];
      40'b?????????????????????????1??????????????:
        _17660_ = b[119:112];
      40'b????????????????????????1???????????????:
        _17660_ = b[127:120];
      40'b???????????????????????1????????????????:
        _17660_ = b[135:128];
      40'b??????????????????????1?????????????????:
        _17660_ = b[143:136];
      40'b?????????????????????1??????????????????:
        _17660_ = b[151:144];
      40'b????????????????????1???????????????????:
        _17660_ = b[159:152];
      40'b???????????????????1????????????????????:
        _17660_ = b[167:160];
      40'b??????????????????1?????????????????????:
        _17660_ = b[175:168];
      40'b?????????????????1??????????????????????:
        _17660_ = b[183:176];
      40'b????????????????1???????????????????????:
        _17660_ = b[191:184];
      40'b???????????????1????????????????????????:
        _17660_ = b[199:192];
      40'b??????????????1?????????????????????????:
        _17660_ = b[207:200];
      40'b?????????????1??????????????????????????:
        _17660_ = b[215:208];
      40'b????????????1???????????????????????????:
        _17660_ = b[223:216];
      40'b???????????1????????????????????????????:
        _17660_ = b[231:224];
      40'b??????????1?????????????????????????????:
        _17660_ = b[239:232];
      40'b?????????1??????????????????????????????:
        _17660_ = b[247:240];
      40'b????????1???????????????????????????????:
        _17660_ = b[255:248];
      40'b???????1????????????????????????????????:
        _17660_ = b[263:256];
      40'b??????1?????????????????????????????????:
        _17660_ = b[271:264];
      40'b?????1??????????????????????????????????:
        _17660_ = b[279:272];
      40'b????1???????????????????????????????????:
        _17660_ = b[287:280];
      40'b???1????????????????????????????????????:
        _17660_ = b[295:288];
      40'b??1?????????????????????????????????????:
        _17660_ = b[303:296];
      40'b?1??????????????????????????????????????:
        _17660_ = b[311:304];
      40'b1???????????????????????????????????????:
        _17660_ = b[319:312];
      default:
        _17660_ = a;
    endcase
  endfunction
  assign vec_data_039 = _17660_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304], data_d1[319:312] }, { _08221_, _08220_, _08219_, _08218_, _08217_, _08216_, _08215_, _08214_, _08213_, _08212_, _08211_, _08210_, _08209_, _08208_, _08207_, _08206_, _08205_, _08204_, _08203_, _08202_, _08201_, _08200_, _08199_, _08198_, _08197_, _08196_, _08195_, _08194_, _08193_, _08192_, _08191_, _08190_, _08189_, _08188_, _08187_, _08186_, _08185_, _08184_, _08183_, _08182_ });
  assign _08182_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5023|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b101000;
  assign _08183_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5022|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100111;
  assign _08184_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5021|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100110;
  assign _08185_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5020|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100101;
  assign _08186_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5019|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100100;
  assign _08187_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100011;
  assign _08188_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100010;
  assign _08189_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100001;
  assign _08190_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 6'b100000;
  assign _08191_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11111;
  assign _08192_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11110;
  assign _08193_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11101;
  assign _08194_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11100;
  assign _08195_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11011;
  assign _08196_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11010;
  assign _08197_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5008|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11001;
  assign _08198_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5007|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b11000;
  assign _08199_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5006|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10111;
  assign _08200_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5005|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10110;
  assign _08201_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5004|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10101;
  assign _08202_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5003|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10100;
  assign _08203_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5002|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10011;
  assign _08204_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5001|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10010;
  assign _08205_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:5000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10001;
  assign _08206_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 5'b10000;
  assign _08207_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1111;
  assign _08208_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1110;
  assign _08209_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1101;
  assign _08210_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1100;
  assign _08211_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1011;
  assign _08212_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1010;
  assign _08213_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1001;
  assign _08214_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4991|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 4'b1000;
  assign _08215_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4990|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 3'b111;
  assign _08216_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4989|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 3'b110;
  assign _08217_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4988|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 3'b101;
  assign _08218_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4987|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 3'b100;
  assign _08219_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4986|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 2'b11;
  assign _08220_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4985|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 2'b10;
  assign _08221_ = vec_sum_039_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4984|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4983" *) 1'b1;
  function [7:0] _17701_;
    input [7:0] a;
    input [311:0] b;
    input [38:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *)
    (* parallel_case *)
    casez (s)
      39'b??????????????????????????????????????1:
        _17701_ = b[7:0];
      39'b?????????????????????????????????????1?:
        _17701_ = b[15:8];
      39'b????????????????????????????????????1??:
        _17701_ = b[23:16];
      39'b???????????????????????????????????1???:
        _17701_ = b[31:24];
      39'b??????????????????????????????????1????:
        _17701_ = b[39:32];
      39'b?????????????????????????????????1?????:
        _17701_ = b[47:40];
      39'b????????????????????????????????1??????:
        _17701_ = b[55:48];
      39'b???????????????????????????????1???????:
        _17701_ = b[63:56];
      39'b??????????????????????????????1????????:
        _17701_ = b[71:64];
      39'b?????????????????????????????1?????????:
        _17701_ = b[79:72];
      39'b????????????????????????????1??????????:
        _17701_ = b[87:80];
      39'b???????????????????????????1???????????:
        _17701_ = b[95:88];
      39'b??????????????????????????1????????????:
        _17701_ = b[103:96];
      39'b?????????????????????????1?????????????:
        _17701_ = b[111:104];
      39'b????????????????????????1??????????????:
        _17701_ = b[119:112];
      39'b???????????????????????1???????????????:
        _17701_ = b[127:120];
      39'b??????????????????????1????????????????:
        _17701_ = b[135:128];
      39'b?????????????????????1?????????????????:
        _17701_ = b[143:136];
      39'b????????????????????1??????????????????:
        _17701_ = b[151:144];
      39'b???????????????????1???????????????????:
        _17701_ = b[159:152];
      39'b??????????????????1????????????????????:
        _17701_ = b[167:160];
      39'b?????????????????1?????????????????????:
        _17701_ = b[175:168];
      39'b????????????????1??????????????????????:
        _17701_ = b[183:176];
      39'b???????????????1???????????????????????:
        _17701_ = b[191:184];
      39'b??????????????1????????????????????????:
        _17701_ = b[199:192];
      39'b?????????????1?????????????????????????:
        _17701_ = b[207:200];
      39'b????????????1??????????????????????????:
        _17701_ = b[215:208];
      39'b???????????1???????????????????????????:
        _17701_ = b[223:216];
      39'b??????????1????????????????????????????:
        _17701_ = b[231:224];
      39'b?????????1?????????????????????????????:
        _17701_ = b[239:232];
      39'b????????1??????????????????????????????:
        _17701_ = b[247:240];
      39'b???????1???????????????????????????????:
        _17701_ = b[255:248];
      39'b??????1????????????????????????????????:
        _17701_ = b[263:256];
      39'b?????1?????????????????????????????????:
        _17701_ = b[271:264];
      39'b????1??????????????????????????????????:
        _17701_ = b[279:272];
      39'b???1???????????????????????????????????:
        _17701_ = b[287:280];
      39'b??1????????????????????????????????????:
        _17701_ = b[295:288];
      39'b?1?????????????????????????????????????:
        _17701_ = b[303:296];
      39'b1??????????????????????????????????????:
        _17701_ = b[311:304];
      default:
        _17701_ = a;
    endcase
  endfunction
  assign vec_data_038 = _17701_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296], data_d1[311:304] }, { _08260_, _08259_, _08258_, _08257_, _08256_, _08255_, _08254_, _08253_, _08252_, _08251_, _08250_, _08249_, _08248_, _08247_, _08246_, _08245_, _08244_, _08243_, _08242_, _08241_, _08240_, _08239_, _08238_, _08237_, _08236_, _08235_, _08234_, _08233_, _08232_, _08231_, _08230_, _08229_, _08228_, _08227_, _08226_, _08225_, _08224_, _08223_, _08222_ });
  assign _08222_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4975|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100111;
  assign _08223_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4974|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100110;
  assign _08224_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4973|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100101;
  assign _08225_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4972|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100100;
  assign _08226_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4971|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100011;
  assign _08227_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4970|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100010;
  assign _08228_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4969|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100001;
  assign _08229_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4968|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 6'b100000;
  assign _08230_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11111;
  assign _08231_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11110;
  assign _08232_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11101;
  assign _08233_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11100;
  assign _08234_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11011;
  assign _08235_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11010;
  assign _08236_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11001;
  assign _08237_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4960|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b11000;
  assign _08238_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4959|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10111;
  assign _08239_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4958|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10110;
  assign _08240_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4957|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10101;
  assign _08241_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4956|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10100;
  assign _08242_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4955|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10011;
  assign _08243_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4954|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10010;
  assign _08244_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4953|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10001;
  assign _08245_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 5'b10000;
  assign _08246_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1111;
  assign _08247_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1110;
  assign _08248_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1101;
  assign _08249_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1100;
  assign _08250_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1011;
  assign _08251_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4946|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1010;
  assign _08252_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4945|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1001;
  assign _08253_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4944|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 4'b1000;
  assign _08254_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4943|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 3'b111;
  assign _08255_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4942|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 3'b110;
  assign _08256_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4941|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 3'b101;
  assign _08257_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4940|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 3'b100;
  assign _08258_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4939|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 2'b11;
  assign _08259_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 2'b10;
  assign _08260_ = vec_sum_038_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4936" *) 1'b1;
  function [7:0] _17741_;
    input [7:0] a;
    input [303:0] b;
    input [37:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *)
    (* parallel_case *)
    casez (s)
      38'b?????????????????????????????????????1:
        _17741_ = b[7:0];
      38'b????????????????????????????????????1?:
        _17741_ = b[15:8];
      38'b???????????????????????????????????1??:
        _17741_ = b[23:16];
      38'b??????????????????????????????????1???:
        _17741_ = b[31:24];
      38'b?????????????????????????????????1????:
        _17741_ = b[39:32];
      38'b????????????????????????????????1?????:
        _17741_ = b[47:40];
      38'b???????????????????????????????1??????:
        _17741_ = b[55:48];
      38'b??????????????????????????????1???????:
        _17741_ = b[63:56];
      38'b?????????????????????????????1????????:
        _17741_ = b[71:64];
      38'b????????????????????????????1?????????:
        _17741_ = b[79:72];
      38'b???????????????????????????1??????????:
        _17741_ = b[87:80];
      38'b??????????????????????????1???????????:
        _17741_ = b[95:88];
      38'b?????????????????????????1????????????:
        _17741_ = b[103:96];
      38'b????????????????????????1?????????????:
        _17741_ = b[111:104];
      38'b???????????????????????1??????????????:
        _17741_ = b[119:112];
      38'b??????????????????????1???????????????:
        _17741_ = b[127:120];
      38'b?????????????????????1????????????????:
        _17741_ = b[135:128];
      38'b????????????????????1?????????????????:
        _17741_ = b[143:136];
      38'b???????????????????1??????????????????:
        _17741_ = b[151:144];
      38'b??????????????????1???????????????????:
        _17741_ = b[159:152];
      38'b?????????????????1????????????????????:
        _17741_ = b[167:160];
      38'b????????????????1?????????????????????:
        _17741_ = b[175:168];
      38'b???????????????1??????????????????????:
        _17741_ = b[183:176];
      38'b??????????????1???????????????????????:
        _17741_ = b[191:184];
      38'b?????????????1????????????????????????:
        _17741_ = b[199:192];
      38'b????????????1?????????????????????????:
        _17741_ = b[207:200];
      38'b???????????1??????????????????????????:
        _17741_ = b[215:208];
      38'b??????????1???????????????????????????:
        _17741_ = b[223:216];
      38'b?????????1????????????????????????????:
        _17741_ = b[231:224];
      38'b????????1?????????????????????????????:
        _17741_ = b[239:232];
      38'b???????1??????????????????????????????:
        _17741_ = b[247:240];
      38'b??????1???????????????????????????????:
        _17741_ = b[255:248];
      38'b?????1????????????????????????????????:
        _17741_ = b[263:256];
      38'b????1?????????????????????????????????:
        _17741_ = b[271:264];
      38'b???1??????????????????????????????????:
        _17741_ = b[279:272];
      38'b??1???????????????????????????????????:
        _17741_ = b[287:280];
      38'b?1????????????????????????????????????:
        _17741_ = b[295:288];
      38'b1?????????????????????????????????????:
        _17741_ = b[303:296];
      default:
        _17741_ = a;
    endcase
  endfunction
  assign vec_data_037 = _17741_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288], data_d1[303:296] }, { _08298_, _08297_, _08296_, _08295_, _08294_, _08293_, _08292_, _08291_, _08290_, _08289_, _08288_, _08287_, _08286_, _08285_, _08284_, _08283_, _08282_, _08281_, _08280_, _08279_, _08278_, _08277_, _08276_, _08275_, _08274_, _08273_, _08272_, _08271_, _08270_, _08269_, _08268_, _08267_, _08266_, _08265_, _08264_, _08263_, _08262_, _08261_ });
  assign _08261_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4928|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100110;
  assign _08262_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4927|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100101;
  assign _08263_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4926|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100100;
  assign _08264_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100011;
  assign _08265_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100010;
  assign _08266_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100001;
  assign _08267_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 6'b100000;
  assign _08268_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4921|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11111;
  assign _08269_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4920|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11110;
  assign _08270_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4919|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11101;
  assign _08271_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4918|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11100;
  assign _08272_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4917|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11011;
  assign _08273_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4916|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11010;
  assign _08274_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4915|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11001;
  assign _08275_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4914|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b11000;
  assign _08276_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10111;
  assign _08277_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10110;
  assign _08278_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10101;
  assign _08279_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4910|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10100;
  assign _08280_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4909|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10011;
  assign _08281_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4908|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10010;
  assign _08282_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4907|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10001;
  assign _08283_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4906|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 5'b10000;
  assign _08284_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4905|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1111;
  assign _08285_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4904|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1110;
  assign _08286_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4903|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1101;
  assign _08287_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1100;
  assign _08288_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1011;
  assign _08289_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4900|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1010;
  assign _08290_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4899|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1001;
  assign _08291_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4898|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 4'b1000;
  assign _08292_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4897|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 3'b111;
  assign _08293_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4896|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 3'b110;
  assign _08294_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4895|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 3'b101;
  assign _08295_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4894|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 3'b100;
  assign _08296_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4893|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 2'b11;
  assign _08297_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 2'b10;
  assign _08298_ = vec_sum_037_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4891|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4890" *) 1'b1;
  function [7:0] _17780_;
    input [7:0] a;
    input [295:0] b;
    input [36:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *)
    (* parallel_case *)
    casez (s)
      37'b????????????????????????????????????1:
        _17780_ = b[7:0];
      37'b???????????????????????????????????1?:
        _17780_ = b[15:8];
      37'b??????????????????????????????????1??:
        _17780_ = b[23:16];
      37'b?????????????????????????????????1???:
        _17780_ = b[31:24];
      37'b????????????????????????????????1????:
        _17780_ = b[39:32];
      37'b???????????????????????????????1?????:
        _17780_ = b[47:40];
      37'b??????????????????????????????1??????:
        _17780_ = b[55:48];
      37'b?????????????????????????????1???????:
        _17780_ = b[63:56];
      37'b????????????????????????????1????????:
        _17780_ = b[71:64];
      37'b???????????????????????????1?????????:
        _17780_ = b[79:72];
      37'b??????????????????????????1??????????:
        _17780_ = b[87:80];
      37'b?????????????????????????1???????????:
        _17780_ = b[95:88];
      37'b????????????????????????1????????????:
        _17780_ = b[103:96];
      37'b???????????????????????1?????????????:
        _17780_ = b[111:104];
      37'b??????????????????????1??????????????:
        _17780_ = b[119:112];
      37'b?????????????????????1???????????????:
        _17780_ = b[127:120];
      37'b????????????????????1????????????????:
        _17780_ = b[135:128];
      37'b???????????????????1?????????????????:
        _17780_ = b[143:136];
      37'b??????????????????1??????????????????:
        _17780_ = b[151:144];
      37'b?????????????????1???????????????????:
        _17780_ = b[159:152];
      37'b????????????????1????????????????????:
        _17780_ = b[167:160];
      37'b???????????????1?????????????????????:
        _17780_ = b[175:168];
      37'b??????????????1??????????????????????:
        _17780_ = b[183:176];
      37'b?????????????1???????????????????????:
        _17780_ = b[191:184];
      37'b????????????1????????????????????????:
        _17780_ = b[199:192];
      37'b???????????1?????????????????????????:
        _17780_ = b[207:200];
      37'b??????????1??????????????????????????:
        _17780_ = b[215:208];
      37'b?????????1???????????????????????????:
        _17780_ = b[223:216];
      37'b????????1????????????????????????????:
        _17780_ = b[231:224];
      37'b???????1?????????????????????????????:
        _17780_ = b[239:232];
      37'b??????1??????????????????????????????:
        _17780_ = b[247:240];
      37'b?????1???????????????????????????????:
        _17780_ = b[255:248];
      37'b????1????????????????????????????????:
        _17780_ = b[263:256];
      37'b???1?????????????????????????????????:
        _17780_ = b[271:264];
      37'b??1??????????????????????????????????:
        _17780_ = b[279:272];
      37'b?1???????????????????????????????????:
        _17780_ = b[287:280];
      37'b1????????????????????????????????????:
        _17780_ = b[295:288];
      default:
        _17780_ = a;
    endcase
  endfunction
  assign vec_data_036 = _17780_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280], data_d1[295:288] }, { _08335_, _08334_, _08333_, _08332_, _08331_, _08330_, _08329_, _08328_, _08327_, _08326_, _08325_, _08324_, _08323_, _08322_, _08321_, _08320_, _08319_, _08318_, _08317_, _08316_, _08315_, _08314_, _08313_, _08312_, _08311_, _08310_, _08309_, _08308_, _08307_, _08306_, _08305_, _08304_, _08303_, _08302_, _08301_, _08300_, _08299_ });
  assign _08299_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4882|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100101;
  assign _08300_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4881|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100100;
  assign _08301_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4880|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100011;
  assign _08302_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4879|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100010;
  assign _08303_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4878|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100001;
  assign _08304_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4877|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 6'b100000;
  assign _08305_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4876|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11111;
  assign _08306_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4875|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11110;
  assign _08307_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4874|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11101;
  assign _08308_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4873|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11100;
  assign _08309_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4872|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11011;
  assign _08310_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4871|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11010;
  assign _08311_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4870|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11001;
  assign _08312_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4869|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b11000;
  assign _08313_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4868|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10111;
  assign _08314_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4867|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10110;
  assign _08315_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4866|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10101;
  assign _08316_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4865|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10100;
  assign _08317_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4864|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10011;
  assign _08318_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4863|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10010;
  assign _08319_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4862|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10001;
  assign _08320_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4861|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 5'b10000;
  assign _08321_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4860|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1111;
  assign _08322_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4859|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1110;
  assign _08323_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4858|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1101;
  assign _08324_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4857|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1100;
  assign _08325_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4856|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1011;
  assign _08326_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4855|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1010;
  assign _08327_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4854|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1001;
  assign _08328_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4853|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 4'b1000;
  assign _08329_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4852|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 3'b111;
  assign _08330_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4851|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 3'b110;
  assign _08331_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4850|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 3'b101;
  assign _08332_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4849|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 3'b100;
  assign _08333_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4848|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 2'b11;
  assign _08334_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4847|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 2'b10;
  assign _08335_ = vec_sum_036_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4846|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4845" *) 1'b1;
  function [7:0] _17818_;
    input [7:0] a;
    input [287:0] b;
    input [35:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *)
    (* parallel_case *)
    casez (s)
      36'b???????????????????????????????????1:
        _17818_ = b[7:0];
      36'b??????????????????????????????????1?:
        _17818_ = b[15:8];
      36'b?????????????????????????????????1??:
        _17818_ = b[23:16];
      36'b????????????????????????????????1???:
        _17818_ = b[31:24];
      36'b???????????????????????????????1????:
        _17818_ = b[39:32];
      36'b??????????????????????????????1?????:
        _17818_ = b[47:40];
      36'b?????????????????????????????1??????:
        _17818_ = b[55:48];
      36'b????????????????????????????1???????:
        _17818_ = b[63:56];
      36'b???????????????????????????1????????:
        _17818_ = b[71:64];
      36'b??????????????????????????1?????????:
        _17818_ = b[79:72];
      36'b?????????????????????????1??????????:
        _17818_ = b[87:80];
      36'b????????????????????????1???????????:
        _17818_ = b[95:88];
      36'b???????????????????????1????????????:
        _17818_ = b[103:96];
      36'b??????????????????????1?????????????:
        _17818_ = b[111:104];
      36'b?????????????????????1??????????????:
        _17818_ = b[119:112];
      36'b????????????????????1???????????????:
        _17818_ = b[127:120];
      36'b???????????????????1????????????????:
        _17818_ = b[135:128];
      36'b??????????????????1?????????????????:
        _17818_ = b[143:136];
      36'b?????????????????1??????????????????:
        _17818_ = b[151:144];
      36'b????????????????1???????????????????:
        _17818_ = b[159:152];
      36'b???????????????1????????????????????:
        _17818_ = b[167:160];
      36'b??????????????1?????????????????????:
        _17818_ = b[175:168];
      36'b?????????????1??????????????????????:
        _17818_ = b[183:176];
      36'b????????????1???????????????????????:
        _17818_ = b[191:184];
      36'b???????????1????????????????????????:
        _17818_ = b[199:192];
      36'b??????????1?????????????????????????:
        _17818_ = b[207:200];
      36'b?????????1??????????????????????????:
        _17818_ = b[215:208];
      36'b????????1???????????????????????????:
        _17818_ = b[223:216];
      36'b???????1????????????????????????????:
        _17818_ = b[231:224];
      36'b??????1?????????????????????????????:
        _17818_ = b[239:232];
      36'b?????1??????????????????????????????:
        _17818_ = b[247:240];
      36'b????1???????????????????????????????:
        _17818_ = b[255:248];
      36'b???1????????????????????????????????:
        _17818_ = b[263:256];
      36'b??1?????????????????????????????????:
        _17818_ = b[271:264];
      36'b?1??????????????????????????????????:
        _17818_ = b[279:272];
      36'b1???????????????????????????????????:
        _17818_ = b[287:280];
      default:
        _17818_ = a;
    endcase
  endfunction
  assign vec_data_035 = _17818_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272], data_d1[287:280] }, { _08371_, _08370_, _08369_, _08368_, _08367_, _08366_, _08365_, _08364_, _08363_, _08362_, _08361_, _08360_, _08359_, _08358_, _08357_, _08356_, _08355_, _08354_, _08353_, _08352_, _08351_, _08350_, _08349_, _08348_, _08347_, _08346_, _08345_, _08344_, _08343_, _08342_, _08341_, _08340_, _08339_, _08338_, _08337_, _08336_ });
  assign _08336_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4837|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 6'b100100;
  assign _08337_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4836|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 6'b100011;
  assign _08338_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4835|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 6'b100010;
  assign _08339_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4834|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 6'b100001;
  assign _08340_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4833|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 6'b100000;
  assign _08341_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4832|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11111;
  assign _08342_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4831|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11110;
  assign _08343_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4830|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11101;
  assign _08344_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4829|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11100;
  assign _08345_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4828|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11011;
  assign _08346_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4827|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11010;
  assign _08347_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4826|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11001;
  assign _08348_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4825|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b11000;
  assign _08349_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4824|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10111;
  assign _08350_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4823|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10110;
  assign _08351_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4822|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10101;
  assign _08352_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4821|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10100;
  assign _08353_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4820|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10011;
  assign _08354_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4819|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10010;
  assign _08355_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4818|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10001;
  assign _08356_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4817|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 5'b10000;
  assign _08357_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4816|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1111;
  assign _08358_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4815|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1110;
  assign _08359_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4814|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1101;
  assign _08360_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4813|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1100;
  assign _08361_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4812|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1011;
  assign _08362_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4811|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1010;
  assign _08363_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4810|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1001;
  assign _08364_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4809|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 4'b1000;
  assign _08365_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4808|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 3'b111;
  assign _08366_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4807|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 3'b110;
  assign _08367_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4806|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 3'b101;
  assign _08368_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4805|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 3'b100;
  assign _08369_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4804|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 2'b11;
  assign _08370_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4803|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 2'b10;
  assign _08371_ = vec_sum_035_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4802|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4801" *) 1'b1;
  function [7:0] _17855_;
    input [7:0] a;
    input [279:0] b;
    input [34:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *)
    (* parallel_case *)
    casez (s)
      35'b??????????????????????????????????1:
        _17855_ = b[7:0];
      35'b?????????????????????????????????1?:
        _17855_ = b[15:8];
      35'b????????????????????????????????1??:
        _17855_ = b[23:16];
      35'b???????????????????????????????1???:
        _17855_ = b[31:24];
      35'b??????????????????????????????1????:
        _17855_ = b[39:32];
      35'b?????????????????????????????1?????:
        _17855_ = b[47:40];
      35'b????????????????????????????1??????:
        _17855_ = b[55:48];
      35'b???????????????????????????1???????:
        _17855_ = b[63:56];
      35'b??????????????????????????1????????:
        _17855_ = b[71:64];
      35'b?????????????????????????1?????????:
        _17855_ = b[79:72];
      35'b????????????????????????1??????????:
        _17855_ = b[87:80];
      35'b???????????????????????1???????????:
        _17855_ = b[95:88];
      35'b??????????????????????1????????????:
        _17855_ = b[103:96];
      35'b?????????????????????1?????????????:
        _17855_ = b[111:104];
      35'b????????????????????1??????????????:
        _17855_ = b[119:112];
      35'b???????????????????1???????????????:
        _17855_ = b[127:120];
      35'b??????????????????1????????????????:
        _17855_ = b[135:128];
      35'b?????????????????1?????????????????:
        _17855_ = b[143:136];
      35'b????????????????1??????????????????:
        _17855_ = b[151:144];
      35'b???????????????1???????????????????:
        _17855_ = b[159:152];
      35'b??????????????1????????????????????:
        _17855_ = b[167:160];
      35'b?????????????1?????????????????????:
        _17855_ = b[175:168];
      35'b????????????1??????????????????????:
        _17855_ = b[183:176];
      35'b???????????1???????????????????????:
        _17855_ = b[191:184];
      35'b??????????1????????????????????????:
        _17855_ = b[199:192];
      35'b?????????1?????????????????????????:
        _17855_ = b[207:200];
      35'b????????1??????????????????????????:
        _17855_ = b[215:208];
      35'b???????1???????????????????????????:
        _17855_ = b[223:216];
      35'b??????1????????????????????????????:
        _17855_ = b[231:224];
      35'b?????1?????????????????????????????:
        _17855_ = b[239:232];
      35'b????1??????????????????????????????:
        _17855_ = b[247:240];
      35'b???1???????????????????????????????:
        _17855_ = b[255:248];
      35'b??1????????????????????????????????:
        _17855_ = b[263:256];
      35'b?1?????????????????????????????????:
        _17855_ = b[271:264];
      35'b1??????????????????????????????????:
        _17855_ = b[279:272];
      default:
        _17855_ = a;
    endcase
  endfunction
  assign vec_data_034 = _17855_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264], data_d1[279:272] }, { _08406_, _08405_, _08404_, _08403_, _08402_, _08401_, _08400_, _08399_, _08398_, _08397_, _08396_, _08395_, _08394_, _08393_, _08392_, _08391_, _08390_, _08389_, _08388_, _08387_, _08386_, _08385_, _08384_, _08383_, _08382_, _08381_, _08380_, _08379_, _08378_, _08377_, _08376_, _08375_, _08374_, _08373_, _08372_ });
  assign _08372_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4793|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 6'b100011;
  assign _08373_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4792|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 6'b100010;
  assign _08374_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4791|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 6'b100001;
  assign _08375_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4790|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 6'b100000;
  assign _08376_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4789|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11111;
  assign _08377_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4788|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11110;
  assign _08378_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4787|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11101;
  assign _08379_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4786|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11100;
  assign _08380_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4785|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11011;
  assign _08381_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4784|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11010;
  assign _08382_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4783|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11001;
  assign _08383_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4782|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b11000;
  assign _08384_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4781|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10111;
  assign _08385_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4780|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10110;
  assign _08386_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4779|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10101;
  assign _08387_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4778|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10100;
  assign _08388_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4777|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10011;
  assign _08389_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4776|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10010;
  assign _08390_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4775|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10001;
  assign _08391_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4774|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 5'b10000;
  assign _08392_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4773|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1111;
  assign _08393_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4772|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1110;
  assign _08394_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4771|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1101;
  assign _08395_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4770|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1100;
  assign _08396_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4769|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1011;
  assign _08397_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4768|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1010;
  assign _08398_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4767|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1001;
  assign _08399_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4766|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 4'b1000;
  assign _08400_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4765|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 3'b111;
  assign _08401_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4764|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 3'b110;
  assign _08402_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4763|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 3'b101;
  assign _08403_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4762|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 3'b100;
  assign _08404_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4761|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 2'b11;
  assign _08405_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4760|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 2'b10;
  assign _08406_ = vec_sum_034_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4759|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4758" *) 1'b1;
  function [7:0] _17891_;
    input [7:0] a;
    input [271:0] b;
    input [33:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *)
    (* parallel_case *)
    casez (s)
      34'b?????????????????????????????????1:
        _17891_ = b[7:0];
      34'b????????????????????????????????1?:
        _17891_ = b[15:8];
      34'b???????????????????????????????1??:
        _17891_ = b[23:16];
      34'b??????????????????????????????1???:
        _17891_ = b[31:24];
      34'b?????????????????????????????1????:
        _17891_ = b[39:32];
      34'b????????????????????????????1?????:
        _17891_ = b[47:40];
      34'b???????????????????????????1??????:
        _17891_ = b[55:48];
      34'b??????????????????????????1???????:
        _17891_ = b[63:56];
      34'b?????????????????????????1????????:
        _17891_ = b[71:64];
      34'b????????????????????????1?????????:
        _17891_ = b[79:72];
      34'b???????????????????????1??????????:
        _17891_ = b[87:80];
      34'b??????????????????????1???????????:
        _17891_ = b[95:88];
      34'b?????????????????????1????????????:
        _17891_ = b[103:96];
      34'b????????????????????1?????????????:
        _17891_ = b[111:104];
      34'b???????????????????1??????????????:
        _17891_ = b[119:112];
      34'b??????????????????1???????????????:
        _17891_ = b[127:120];
      34'b?????????????????1????????????????:
        _17891_ = b[135:128];
      34'b????????????????1?????????????????:
        _17891_ = b[143:136];
      34'b???????????????1??????????????????:
        _17891_ = b[151:144];
      34'b??????????????1???????????????????:
        _17891_ = b[159:152];
      34'b?????????????1????????????????????:
        _17891_ = b[167:160];
      34'b????????????1?????????????????????:
        _17891_ = b[175:168];
      34'b???????????1??????????????????????:
        _17891_ = b[183:176];
      34'b??????????1???????????????????????:
        _17891_ = b[191:184];
      34'b?????????1????????????????????????:
        _17891_ = b[199:192];
      34'b????????1?????????????????????????:
        _17891_ = b[207:200];
      34'b???????1??????????????????????????:
        _17891_ = b[215:208];
      34'b??????1???????????????????????????:
        _17891_ = b[223:216];
      34'b?????1????????????????????????????:
        _17891_ = b[231:224];
      34'b????1?????????????????????????????:
        _17891_ = b[239:232];
      34'b???1??????????????????????????????:
        _17891_ = b[247:240];
      34'b??1???????????????????????????????:
        _17891_ = b[255:248];
      34'b?1????????????????????????????????:
        _17891_ = b[263:256];
      34'b1?????????????????????????????????:
        _17891_ = b[271:264];
      default:
        _17891_ = a;
    endcase
  endfunction
  assign vec_data_033 = _17891_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256], data_d1[271:264] }, { _08440_, _08439_, _08438_, _08437_, _08436_, _08435_, _08434_, _08433_, _08432_, _08431_, _08430_, _08429_, _08428_, _08427_, _08426_, _08425_, _08424_, _08423_, _08422_, _08421_, _08420_, _08419_, _08418_, _08417_, _08416_, _08415_, _08414_, _08413_, _08412_, _08411_, _08410_, _08409_, _08408_, _08407_ });
  assign _08407_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4750|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 6'b100010;
  assign _08408_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4749|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 6'b100001;
  assign _08409_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4748|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 6'b100000;
  assign _08410_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4747|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11111;
  assign _08411_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4746|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11110;
  assign _08412_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4745|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11101;
  assign _08413_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4744|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11100;
  assign _08414_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4743|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11011;
  assign _08415_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4742|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11010;
  assign _08416_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4741|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11001;
  assign _08417_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4740|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b11000;
  assign _08418_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4739|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10111;
  assign _08419_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4738|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10110;
  assign _08420_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4737|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10101;
  assign _08421_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4736|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10100;
  assign _08422_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4735|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10011;
  assign _08423_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4734|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10010;
  assign _08424_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4733|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10001;
  assign _08425_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4732|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 5'b10000;
  assign _08426_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4731|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1111;
  assign _08427_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4730|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1110;
  assign _08428_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4729|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1101;
  assign _08429_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4728|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1100;
  assign _08430_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4727|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1011;
  assign _08431_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4726|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1010;
  assign _08432_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4725|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1001;
  assign _08433_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4724|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 4'b1000;
  assign _08434_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4723|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 3'b111;
  assign _08435_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4722|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 3'b110;
  assign _08436_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4721|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 3'b101;
  assign _08437_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4720|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 3'b100;
  assign _08438_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4719|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 2'b11;
  assign _08439_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4718|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 2'b10;
  assign _08440_ = vec_sum_033_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4717|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4716" *) 1'b1;
  function [7:0] _17926_;
    input [7:0] a;
    input [263:0] b;
    input [32:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *)
    (* parallel_case *)
    casez (s)
      33'b????????????????????????????????1:
        _17926_ = b[7:0];
      33'b???????????????????????????????1?:
        _17926_ = b[15:8];
      33'b??????????????????????????????1??:
        _17926_ = b[23:16];
      33'b?????????????????????????????1???:
        _17926_ = b[31:24];
      33'b????????????????????????????1????:
        _17926_ = b[39:32];
      33'b???????????????????????????1?????:
        _17926_ = b[47:40];
      33'b??????????????????????????1??????:
        _17926_ = b[55:48];
      33'b?????????????????????????1???????:
        _17926_ = b[63:56];
      33'b????????????????????????1????????:
        _17926_ = b[71:64];
      33'b???????????????????????1?????????:
        _17926_ = b[79:72];
      33'b??????????????????????1??????????:
        _17926_ = b[87:80];
      33'b?????????????????????1???????????:
        _17926_ = b[95:88];
      33'b????????????????????1????????????:
        _17926_ = b[103:96];
      33'b???????????????????1?????????????:
        _17926_ = b[111:104];
      33'b??????????????????1??????????????:
        _17926_ = b[119:112];
      33'b?????????????????1???????????????:
        _17926_ = b[127:120];
      33'b????????????????1????????????????:
        _17926_ = b[135:128];
      33'b???????????????1?????????????????:
        _17926_ = b[143:136];
      33'b??????????????1??????????????????:
        _17926_ = b[151:144];
      33'b?????????????1???????????????????:
        _17926_ = b[159:152];
      33'b????????????1????????????????????:
        _17926_ = b[167:160];
      33'b???????????1?????????????????????:
        _17926_ = b[175:168];
      33'b??????????1??????????????????????:
        _17926_ = b[183:176];
      33'b?????????1???????????????????????:
        _17926_ = b[191:184];
      33'b????????1????????????????????????:
        _17926_ = b[199:192];
      33'b???????1?????????????????????????:
        _17926_ = b[207:200];
      33'b??????1??????????????????????????:
        _17926_ = b[215:208];
      33'b?????1???????????????????????????:
        _17926_ = b[223:216];
      33'b????1????????????????????????????:
        _17926_ = b[231:224];
      33'b???1?????????????????????????????:
        _17926_ = b[239:232];
      33'b??1??????????????????????????????:
        _17926_ = b[247:240];
      33'b?1???????????????????????????????:
        _17926_ = b[255:248];
      33'b1????????????????????????????????:
        _17926_ = b[263:256];
      default:
        _17926_ = a;
    endcase
  endfunction
  assign vec_data_032 = _17926_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248], data_d1[263:256] }, { _08473_, _08472_, _08471_, _08470_, _08469_, _08468_, _08467_, _08466_, _08465_, _08464_, _08463_, _08462_, _08461_, _08460_, _08459_, _08458_, _08457_, _08456_, _08455_, _08454_, _08453_, _08452_, _08451_, _08450_, _08449_, _08448_, _08447_, _08446_, _08445_, _08444_, _08443_, _08442_, _08441_ });
  assign _08441_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4708|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 6'b100001;
  assign _08442_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4707|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 6'b100000;
  assign _08443_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4706|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11111;
  assign _08444_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4705|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11110;
  assign _08445_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4704|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11101;
  assign _08446_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4703|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11100;
  assign _08447_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4702|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11011;
  assign _08448_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4701|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11010;
  assign _08449_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4700|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11001;
  assign _08450_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4699|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b11000;
  assign _08451_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4698|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10111;
  assign _08452_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4697|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10110;
  assign _08453_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4696|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10101;
  assign _08454_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4695|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10100;
  assign _08455_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4694|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10011;
  assign _08456_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4693|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10010;
  assign _08457_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4692|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10001;
  assign _08458_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4691|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 5'b10000;
  assign _08459_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4690|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1111;
  assign _08460_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4689|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1110;
  assign _08461_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4688|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1101;
  assign _08462_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4687|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1100;
  assign _08463_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4686|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1011;
  assign _08464_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4685|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1010;
  assign _08465_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4684|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1001;
  assign _08466_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4683|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 4'b1000;
  assign _08467_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4682|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 3'b111;
  assign _08468_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4681|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 3'b110;
  assign _08469_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4680|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 3'b101;
  assign _08470_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4679|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 3'b100;
  assign _08471_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4678|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 2'b11;
  assign _08472_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4677|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 2'b10;
  assign _08473_ = vec_sum_032_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4676|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4675" *) 1'b1;
  function [7:0] _17960_;
    input [7:0] a;
    input [255:0] b;
    input [31:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *)
    (* parallel_case *)
    casez (s)
      32'b???????????????????????????????1:
        _17960_ = b[7:0];
      32'b??????????????????????????????1?:
        _17960_ = b[15:8];
      32'b?????????????????????????????1??:
        _17960_ = b[23:16];
      32'b????????????????????????????1???:
        _17960_ = b[31:24];
      32'b???????????????????????????1????:
        _17960_ = b[39:32];
      32'b??????????????????????????1?????:
        _17960_ = b[47:40];
      32'b?????????????????????????1??????:
        _17960_ = b[55:48];
      32'b????????????????????????1???????:
        _17960_ = b[63:56];
      32'b???????????????????????1????????:
        _17960_ = b[71:64];
      32'b??????????????????????1?????????:
        _17960_ = b[79:72];
      32'b?????????????????????1??????????:
        _17960_ = b[87:80];
      32'b????????????????????1???????????:
        _17960_ = b[95:88];
      32'b???????????????????1????????????:
        _17960_ = b[103:96];
      32'b??????????????????1?????????????:
        _17960_ = b[111:104];
      32'b?????????????????1??????????????:
        _17960_ = b[119:112];
      32'b????????????????1???????????????:
        _17960_ = b[127:120];
      32'b???????????????1????????????????:
        _17960_ = b[135:128];
      32'b??????????????1?????????????????:
        _17960_ = b[143:136];
      32'b?????????????1??????????????????:
        _17960_ = b[151:144];
      32'b????????????1???????????????????:
        _17960_ = b[159:152];
      32'b???????????1????????????????????:
        _17960_ = b[167:160];
      32'b??????????1?????????????????????:
        _17960_ = b[175:168];
      32'b?????????1??????????????????????:
        _17960_ = b[183:176];
      32'b????????1???????????????????????:
        _17960_ = b[191:184];
      32'b???????1????????????????????????:
        _17960_ = b[199:192];
      32'b??????1?????????????????????????:
        _17960_ = b[207:200];
      32'b?????1??????????????????????????:
        _17960_ = b[215:208];
      32'b????1???????????????????????????:
        _17960_ = b[223:216];
      32'b???1????????????????????????????:
        _17960_ = b[231:224];
      32'b??1?????????????????????????????:
        _17960_ = b[239:232];
      32'b?1??????????????????????????????:
        _17960_ = b[247:240];
      32'b1???????????????????????????????:
        _17960_ = b[255:248];
      default:
        _17960_ = a;
    endcase
  endfunction
  assign vec_data_031 = _17960_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240], data_d1[255:248] }, { _08505_, _08504_, _08503_, _08502_, _08501_, _08500_, _08499_, _08498_, _08497_, _08496_, _08495_, _08494_, _08493_, _08492_, _08491_, _08490_, _08489_, _08488_, _08487_, _08486_, _08485_, _08484_, _08483_, _08482_, _08481_, _08480_, _08479_, _08478_, _08477_, _08476_, _08475_, _08474_ });
  assign _08474_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4667|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 6'b100000;
  assign _08475_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4666|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11111;
  assign _08476_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4665|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11110;
  assign _08477_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4664|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11101;
  assign _08478_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4663|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11100;
  assign _08479_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4662|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11011;
  assign _08480_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4661|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11010;
  assign _08481_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4660|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11001;
  assign _08482_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4659|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b11000;
  assign _08483_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4658|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10111;
  assign _08484_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4657|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10110;
  assign _08485_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4656|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10101;
  assign _08486_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4655|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10100;
  assign _08487_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4654|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10011;
  assign _08488_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4653|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10010;
  assign _08489_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4652|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10001;
  assign _08490_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4651|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 5'b10000;
  assign _08491_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4650|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1111;
  assign _08492_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4649|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1110;
  assign _08493_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4648|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1101;
  assign _08494_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4647|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1100;
  assign _08495_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4646|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1011;
  assign _08496_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4645|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1010;
  assign _08497_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4644|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1001;
  assign _08498_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4643|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 4'b1000;
  assign _08499_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4642|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 3'b111;
  assign _08500_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4641|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 3'b110;
  assign _08501_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4640|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 3'b101;
  assign _08502_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4639|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 3'b100;
  assign _08503_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4638|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 2'b11;
  assign _08504_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4637|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 2'b10;
  assign _08505_ = vec_sum_031_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4636|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4635" *) 1'b1;
  function [7:0] _17993_;
    input [7:0] a;
    input [247:0] b;
    input [30:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *)
    (* parallel_case *)
    casez (s)
      31'b??????????????????????????????1:
        _17993_ = b[7:0];
      31'b?????????????????????????????1?:
        _17993_ = b[15:8];
      31'b????????????????????????????1??:
        _17993_ = b[23:16];
      31'b???????????????????????????1???:
        _17993_ = b[31:24];
      31'b??????????????????????????1????:
        _17993_ = b[39:32];
      31'b?????????????????????????1?????:
        _17993_ = b[47:40];
      31'b????????????????????????1??????:
        _17993_ = b[55:48];
      31'b???????????????????????1???????:
        _17993_ = b[63:56];
      31'b??????????????????????1????????:
        _17993_ = b[71:64];
      31'b?????????????????????1?????????:
        _17993_ = b[79:72];
      31'b????????????????????1??????????:
        _17993_ = b[87:80];
      31'b???????????????????1???????????:
        _17993_ = b[95:88];
      31'b??????????????????1????????????:
        _17993_ = b[103:96];
      31'b?????????????????1?????????????:
        _17993_ = b[111:104];
      31'b????????????????1??????????????:
        _17993_ = b[119:112];
      31'b???????????????1???????????????:
        _17993_ = b[127:120];
      31'b??????????????1????????????????:
        _17993_ = b[135:128];
      31'b?????????????1?????????????????:
        _17993_ = b[143:136];
      31'b????????????1??????????????????:
        _17993_ = b[151:144];
      31'b???????????1???????????????????:
        _17993_ = b[159:152];
      31'b??????????1????????????????????:
        _17993_ = b[167:160];
      31'b?????????1?????????????????????:
        _17993_ = b[175:168];
      31'b????????1??????????????????????:
        _17993_ = b[183:176];
      31'b???????1???????????????????????:
        _17993_ = b[191:184];
      31'b??????1????????????????????????:
        _17993_ = b[199:192];
      31'b?????1?????????????????????????:
        _17993_ = b[207:200];
      31'b????1??????????????????????????:
        _17993_ = b[215:208];
      31'b???1???????????????????????????:
        _17993_ = b[223:216];
      31'b??1????????????????????????????:
        _17993_ = b[231:224];
      31'b?1?????????????????????????????:
        _17993_ = b[239:232];
      31'b1??????????????????????????????:
        _17993_ = b[247:240];
      default:
        _17993_ = a;
    endcase
  endfunction
  assign vec_data_030 = _17993_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232], data_d1[247:240] }, { _08536_, _08535_, _08534_, _08533_, _08532_, _08531_, _08530_, _08529_, _08528_, _08527_, _08526_, _08525_, _08524_, _08523_, _08522_, _08521_, _08520_, _08519_, _08518_, _08517_, _08516_, _08515_, _08514_, _08513_, _08512_, _08511_, _08510_, _08509_, _08508_, _08507_, _08506_ });
  assign _08506_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4627|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11111;
  assign _08507_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4626|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11110;
  assign _08508_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4625|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11101;
  assign _08509_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4624|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11100;
  assign _08510_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4623|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11011;
  assign _08511_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4622|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11010;
  assign _08512_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4621|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11001;
  assign _08513_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4620|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b11000;
  assign _08514_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4619|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10111;
  assign _08515_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4618|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10110;
  assign _08516_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4617|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10101;
  assign _08517_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4616|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10100;
  assign _08518_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4615|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10011;
  assign _08519_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4614|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10010;
  assign _08520_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4613|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10001;
  assign _08521_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4612|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 5'b10000;
  assign _08522_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4611|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1111;
  assign _08523_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4610|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1110;
  assign _08524_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4609|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1101;
  assign _08525_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4608|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1100;
  assign _08526_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4607|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1011;
  assign _08527_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4606|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1010;
  assign _08528_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4605|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1001;
  assign _08529_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4604|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 4'b1000;
  assign _08530_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4603|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 3'b111;
  assign _08531_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4602|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 3'b110;
  assign _08532_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4601|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 3'b101;
  assign _08533_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4600|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 3'b100;
  assign _08534_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4599|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 2'b11;
  assign _08535_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4598|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 2'b10;
  assign _08536_ = vec_sum_030_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4597|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4596" *) 1'b1;
  function [7:0] _18025_;
    input [7:0] a;
    input [239:0] b;
    input [29:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *)
    (* parallel_case *)
    casez (s)
      30'b?????????????????????????????1:
        _18025_ = b[7:0];
      30'b????????????????????????????1?:
        _18025_ = b[15:8];
      30'b???????????????????????????1??:
        _18025_ = b[23:16];
      30'b??????????????????????????1???:
        _18025_ = b[31:24];
      30'b?????????????????????????1????:
        _18025_ = b[39:32];
      30'b????????????????????????1?????:
        _18025_ = b[47:40];
      30'b???????????????????????1??????:
        _18025_ = b[55:48];
      30'b??????????????????????1???????:
        _18025_ = b[63:56];
      30'b?????????????????????1????????:
        _18025_ = b[71:64];
      30'b????????????????????1?????????:
        _18025_ = b[79:72];
      30'b???????????????????1??????????:
        _18025_ = b[87:80];
      30'b??????????????????1???????????:
        _18025_ = b[95:88];
      30'b?????????????????1????????????:
        _18025_ = b[103:96];
      30'b????????????????1?????????????:
        _18025_ = b[111:104];
      30'b???????????????1??????????????:
        _18025_ = b[119:112];
      30'b??????????????1???????????????:
        _18025_ = b[127:120];
      30'b?????????????1????????????????:
        _18025_ = b[135:128];
      30'b????????????1?????????????????:
        _18025_ = b[143:136];
      30'b???????????1??????????????????:
        _18025_ = b[151:144];
      30'b??????????1???????????????????:
        _18025_ = b[159:152];
      30'b?????????1????????????????????:
        _18025_ = b[167:160];
      30'b????????1?????????????????????:
        _18025_ = b[175:168];
      30'b???????1??????????????????????:
        _18025_ = b[183:176];
      30'b??????1???????????????????????:
        _18025_ = b[191:184];
      30'b?????1????????????????????????:
        _18025_ = b[199:192];
      30'b????1?????????????????????????:
        _18025_ = b[207:200];
      30'b???1??????????????????????????:
        _18025_ = b[215:208];
      30'b??1???????????????????????????:
        _18025_ = b[223:216];
      30'b?1????????????????????????????:
        _18025_ = b[231:224];
      30'b1?????????????????????????????:
        _18025_ = b[239:232];
      default:
        _18025_ = a;
    endcase
  endfunction
  assign vec_data_029 = _18025_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224], data_d1[239:232] }, { _08566_, _08565_, _08564_, _08563_, _08562_, _08561_, _08560_, _08559_, _08558_, _08557_, _08556_, _08555_, _08554_, _08553_, _08552_, _08551_, _08550_, _08549_, _08548_, _08547_, _08546_, _08545_, _08544_, _08543_, _08542_, _08541_, _08540_, _08539_, _08538_, _08537_ });
  assign _08537_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4588|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11110;
  assign _08538_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4587|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11101;
  assign _08539_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4586|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11100;
  assign _08540_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4585|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11011;
  assign _08541_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4584|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11010;
  assign _08542_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4583|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11001;
  assign _08543_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4582|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b11000;
  assign _08544_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4581|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10111;
  assign _08545_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4580|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10110;
  assign _08546_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4579|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10101;
  assign _08547_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4578|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10100;
  assign _08548_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4577|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10011;
  assign _08549_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4576|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10010;
  assign _08550_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4575|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10001;
  assign _08551_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4574|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 5'b10000;
  assign _08552_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4573|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1111;
  assign _08553_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4572|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1110;
  assign _08554_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4571|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1101;
  assign _08555_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4570|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1100;
  assign _08556_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4569|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1011;
  assign _08557_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4568|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1010;
  assign _08558_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4567|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1001;
  assign _08559_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4566|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 4'b1000;
  assign _08560_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4565|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 3'b111;
  assign _08561_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4564|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 3'b110;
  assign _08562_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4563|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 3'b101;
  assign _08563_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4562|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 3'b100;
  assign _08564_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4561|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 2'b11;
  assign _08565_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4560|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 2'b10;
  assign _08566_ = vec_sum_029_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4559|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4558" *) 1'b1;
  function [7:0] _18056_;
    input [7:0] a;
    input [231:0] b;
    input [28:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *)
    (* parallel_case *)
    casez (s)
      29'b????????????????????????????1:
        _18056_ = b[7:0];
      29'b???????????????????????????1?:
        _18056_ = b[15:8];
      29'b??????????????????????????1??:
        _18056_ = b[23:16];
      29'b?????????????????????????1???:
        _18056_ = b[31:24];
      29'b????????????????????????1????:
        _18056_ = b[39:32];
      29'b???????????????????????1?????:
        _18056_ = b[47:40];
      29'b??????????????????????1??????:
        _18056_ = b[55:48];
      29'b?????????????????????1???????:
        _18056_ = b[63:56];
      29'b????????????????????1????????:
        _18056_ = b[71:64];
      29'b???????????????????1?????????:
        _18056_ = b[79:72];
      29'b??????????????????1??????????:
        _18056_ = b[87:80];
      29'b?????????????????1???????????:
        _18056_ = b[95:88];
      29'b????????????????1????????????:
        _18056_ = b[103:96];
      29'b???????????????1?????????????:
        _18056_ = b[111:104];
      29'b??????????????1??????????????:
        _18056_ = b[119:112];
      29'b?????????????1???????????????:
        _18056_ = b[127:120];
      29'b????????????1????????????????:
        _18056_ = b[135:128];
      29'b???????????1?????????????????:
        _18056_ = b[143:136];
      29'b??????????1??????????????????:
        _18056_ = b[151:144];
      29'b?????????1???????????????????:
        _18056_ = b[159:152];
      29'b????????1????????????????????:
        _18056_ = b[167:160];
      29'b???????1?????????????????????:
        _18056_ = b[175:168];
      29'b??????1??????????????????????:
        _18056_ = b[183:176];
      29'b?????1???????????????????????:
        _18056_ = b[191:184];
      29'b????1????????????????????????:
        _18056_ = b[199:192];
      29'b???1?????????????????????????:
        _18056_ = b[207:200];
      29'b??1??????????????????????????:
        _18056_ = b[215:208];
      29'b?1???????????????????????????:
        _18056_ = b[223:216];
      29'b1????????????????????????????:
        _18056_ = b[231:224];
      default:
        _18056_ = a;
    endcase
  endfunction
  assign vec_data_028 = _18056_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216], data_d1[231:224] }, { _08595_, _08594_, _08593_, _08592_, _08591_, _08590_, _08589_, _08588_, _08587_, _08586_, _08585_, _08584_, _08583_, _08582_, _08581_, _08580_, _08579_, _08578_, _08577_, _08576_, _08575_, _08574_, _08573_, _08572_, _08571_, _08570_, _08569_, _08568_, _08567_ });
  assign _08567_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4550|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11101;
  assign _08568_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4549|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11100;
  assign _08569_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4548|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11011;
  assign _08570_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4547|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11010;
  assign _08571_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4546|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11001;
  assign _08572_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4545|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b11000;
  assign _08573_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4544|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10111;
  assign _08574_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4543|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10110;
  assign _08575_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4542|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10101;
  assign _08576_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4541|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10100;
  assign _08577_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4540|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10011;
  assign _08578_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4539|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10010;
  assign _08579_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4538|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10001;
  assign _08580_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4537|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 5'b10000;
  assign _08581_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4536|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1111;
  assign _08582_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4535|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1110;
  assign _08583_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4534|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1101;
  assign _08584_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4533|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1100;
  assign _08585_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4532|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1011;
  assign _08586_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4531|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1010;
  assign _08587_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4530|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1001;
  assign _08588_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4529|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 4'b1000;
  assign _08589_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4528|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 3'b111;
  assign _08590_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4527|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 3'b110;
  assign _08591_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4526|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 3'b101;
  assign _08592_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4525|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 3'b100;
  assign _08593_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4524|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 2'b11;
  assign _08594_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4523|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 2'b10;
  assign _08595_ = vec_sum_028_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4522|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4521" *) 1'b1;
  function [7:0] _18086_;
    input [7:0] a;
    input [223:0] b;
    input [27:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *)
    (* parallel_case *)
    casez (s)
      28'b???????????????????????????1:
        _18086_ = b[7:0];
      28'b??????????????????????????1?:
        _18086_ = b[15:8];
      28'b?????????????????????????1??:
        _18086_ = b[23:16];
      28'b????????????????????????1???:
        _18086_ = b[31:24];
      28'b???????????????????????1????:
        _18086_ = b[39:32];
      28'b??????????????????????1?????:
        _18086_ = b[47:40];
      28'b?????????????????????1??????:
        _18086_ = b[55:48];
      28'b????????????????????1???????:
        _18086_ = b[63:56];
      28'b???????????????????1????????:
        _18086_ = b[71:64];
      28'b??????????????????1?????????:
        _18086_ = b[79:72];
      28'b?????????????????1??????????:
        _18086_ = b[87:80];
      28'b????????????????1???????????:
        _18086_ = b[95:88];
      28'b???????????????1????????????:
        _18086_ = b[103:96];
      28'b??????????????1?????????????:
        _18086_ = b[111:104];
      28'b?????????????1??????????????:
        _18086_ = b[119:112];
      28'b????????????1???????????????:
        _18086_ = b[127:120];
      28'b???????????1????????????????:
        _18086_ = b[135:128];
      28'b??????????1?????????????????:
        _18086_ = b[143:136];
      28'b?????????1??????????????????:
        _18086_ = b[151:144];
      28'b????????1???????????????????:
        _18086_ = b[159:152];
      28'b???????1????????????????????:
        _18086_ = b[167:160];
      28'b??????1?????????????????????:
        _18086_ = b[175:168];
      28'b?????1??????????????????????:
        _18086_ = b[183:176];
      28'b????1???????????????????????:
        _18086_ = b[191:184];
      28'b???1????????????????????????:
        _18086_ = b[199:192];
      28'b??1?????????????????????????:
        _18086_ = b[207:200];
      28'b?1??????????????????????????:
        _18086_ = b[215:208];
      28'b1???????????????????????????:
        _18086_ = b[223:216];
      default:
        _18086_ = a;
    endcase
  endfunction
  assign vec_data_027 = _18086_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208], data_d1[223:216] }, { _08623_, _08622_, _08621_, _08620_, _08619_, _08618_, _08617_, _08616_, _08615_, _08614_, _08613_, _08612_, _08611_, _08610_, _08609_, _08608_, _08607_, _08606_, _08605_, _08604_, _08603_, _08602_, _08601_, _08600_, _08599_, _08598_, _08597_, _08596_ });
  assign _08596_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4513|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b11100;
  assign _08597_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4512|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b11011;
  assign _08598_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4511|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b11010;
  assign _08599_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4510|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b11001;
  assign _08600_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4509|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b11000;
  assign _08601_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4508|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10111;
  assign _08602_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4507|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10110;
  assign _08603_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4506|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10101;
  assign _08604_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4505|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10100;
  assign _08605_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4504|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10011;
  assign _08606_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4503|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10010;
  assign _08607_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4502|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10001;
  assign _08608_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4501|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 5'b10000;
  assign _08609_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4500|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1111;
  assign _08610_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4499|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1110;
  assign _08611_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4498|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1101;
  assign _08612_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4497|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1100;
  assign _08613_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4496|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1011;
  assign _08614_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4495|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1010;
  assign _08615_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4494|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1001;
  assign _08616_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4493|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 4'b1000;
  assign _08617_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4492|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 3'b111;
  assign _08618_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4491|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 3'b110;
  assign _08619_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4490|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 3'b101;
  assign _08620_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4489|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 3'b100;
  assign _08621_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4488|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 2'b11;
  assign _08622_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4487|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 2'b10;
  assign _08623_ = vec_sum_027_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4486|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4485" *) 1'b1;
  function [7:0] _18115_;
    input [7:0] a;
    input [215:0] b;
    input [26:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *)
    (* parallel_case *)
    casez (s)
      27'b??????????????????????????1:
        _18115_ = b[7:0];
      27'b?????????????????????????1?:
        _18115_ = b[15:8];
      27'b????????????????????????1??:
        _18115_ = b[23:16];
      27'b???????????????????????1???:
        _18115_ = b[31:24];
      27'b??????????????????????1????:
        _18115_ = b[39:32];
      27'b?????????????????????1?????:
        _18115_ = b[47:40];
      27'b????????????????????1??????:
        _18115_ = b[55:48];
      27'b???????????????????1???????:
        _18115_ = b[63:56];
      27'b??????????????????1????????:
        _18115_ = b[71:64];
      27'b?????????????????1?????????:
        _18115_ = b[79:72];
      27'b????????????????1??????????:
        _18115_ = b[87:80];
      27'b???????????????1???????????:
        _18115_ = b[95:88];
      27'b??????????????1????????????:
        _18115_ = b[103:96];
      27'b?????????????1?????????????:
        _18115_ = b[111:104];
      27'b????????????1??????????????:
        _18115_ = b[119:112];
      27'b???????????1???????????????:
        _18115_ = b[127:120];
      27'b??????????1????????????????:
        _18115_ = b[135:128];
      27'b?????????1?????????????????:
        _18115_ = b[143:136];
      27'b????????1??????????????????:
        _18115_ = b[151:144];
      27'b???????1???????????????????:
        _18115_ = b[159:152];
      27'b??????1????????????????????:
        _18115_ = b[167:160];
      27'b?????1?????????????????????:
        _18115_ = b[175:168];
      27'b????1??????????????????????:
        _18115_ = b[183:176];
      27'b???1???????????????????????:
        _18115_ = b[191:184];
      27'b??1????????????????????????:
        _18115_ = b[199:192];
      27'b?1?????????????????????????:
        _18115_ = b[207:200];
      27'b1??????????????????????????:
        _18115_ = b[215:208];
      default:
        _18115_ = a;
    endcase
  endfunction
  assign vec_data_026 = _18115_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200], data_d1[215:208] }, { _08650_, _08649_, _08648_, _08647_, _08646_, _08645_, _08644_, _08643_, _08642_, _08641_, _08640_, _08639_, _08638_, _08637_, _08636_, _08635_, _08634_, _08633_, _08632_, _08631_, _08630_, _08629_, _08628_, _08627_, _08626_, _08625_, _08624_ });
  assign _08624_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4477|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b11011;
  assign _08625_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4476|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b11010;
  assign _08626_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4475|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b11001;
  assign _08627_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4474|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b11000;
  assign _08628_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4473|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10111;
  assign _08629_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4472|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10110;
  assign _08630_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4471|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10101;
  assign _08631_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4470|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10100;
  assign _08632_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4469|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10011;
  assign _08633_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4468|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10010;
  assign _08634_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4467|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10001;
  assign _08635_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4466|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 5'b10000;
  assign _08636_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4465|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1111;
  assign _08637_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4464|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1110;
  assign _08638_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4463|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1101;
  assign _08639_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4462|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1100;
  assign _08640_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4461|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1011;
  assign _08641_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4460|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1010;
  assign _08642_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4459|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1001;
  assign _08643_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4458|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 4'b1000;
  assign _08644_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4457|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 3'b111;
  assign _08645_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4456|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 3'b110;
  assign _08646_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4455|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 3'b101;
  assign _08647_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4454|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 3'b100;
  assign _08648_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4453|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 2'b11;
  assign _08649_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4452|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 2'b10;
  assign _08650_ = vec_sum_026_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4451|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4450" *) 1'b1;
  function [7:0] _18143_;
    input [7:0] a;
    input [207:0] b;
    input [25:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *)
    (* parallel_case *)
    casez (s)
      26'b?????????????????????????1:
        _18143_ = b[7:0];
      26'b????????????????????????1?:
        _18143_ = b[15:8];
      26'b???????????????????????1??:
        _18143_ = b[23:16];
      26'b??????????????????????1???:
        _18143_ = b[31:24];
      26'b?????????????????????1????:
        _18143_ = b[39:32];
      26'b????????????????????1?????:
        _18143_ = b[47:40];
      26'b???????????????????1??????:
        _18143_ = b[55:48];
      26'b??????????????????1???????:
        _18143_ = b[63:56];
      26'b?????????????????1????????:
        _18143_ = b[71:64];
      26'b????????????????1?????????:
        _18143_ = b[79:72];
      26'b???????????????1??????????:
        _18143_ = b[87:80];
      26'b??????????????1???????????:
        _18143_ = b[95:88];
      26'b?????????????1????????????:
        _18143_ = b[103:96];
      26'b????????????1?????????????:
        _18143_ = b[111:104];
      26'b???????????1??????????????:
        _18143_ = b[119:112];
      26'b??????????1???????????????:
        _18143_ = b[127:120];
      26'b?????????1????????????????:
        _18143_ = b[135:128];
      26'b????????1?????????????????:
        _18143_ = b[143:136];
      26'b???????1??????????????????:
        _18143_ = b[151:144];
      26'b??????1???????????????????:
        _18143_ = b[159:152];
      26'b?????1????????????????????:
        _18143_ = b[167:160];
      26'b????1?????????????????????:
        _18143_ = b[175:168];
      26'b???1??????????????????????:
        _18143_ = b[183:176];
      26'b??1???????????????????????:
        _18143_ = b[191:184];
      26'b?1????????????????????????:
        _18143_ = b[199:192];
      26'b1?????????????????????????:
        _18143_ = b[207:200];
      default:
        _18143_ = a;
    endcase
  endfunction
  assign vec_data_025 = _18143_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192], data_d1[207:200] }, { _08676_, _08675_, _08674_, _08673_, _08672_, _08671_, _08670_, _08669_, _08668_, _08667_, _08666_, _08665_, _08664_, _08663_, _08662_, _08661_, _08660_, _08659_, _08658_, _08657_, _08656_, _08655_, _08654_, _08653_, _08652_, _08651_ });
  assign _08651_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4442|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b11010;
  assign _08652_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4441|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b11001;
  assign _08653_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4440|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b11000;
  assign _08654_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4439|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10111;
  assign _08655_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4438|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10110;
  assign _08656_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4437|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10101;
  assign _08657_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4436|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10100;
  assign _08658_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4435|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10011;
  assign _08659_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4434|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10010;
  assign _08660_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4433|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10001;
  assign _08661_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4432|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 5'b10000;
  assign _08662_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4431|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1111;
  assign _08663_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4430|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1110;
  assign _08664_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4429|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1101;
  assign _08665_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4428|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1100;
  assign _08666_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4427|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1011;
  assign _08667_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4426|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1010;
  assign _08668_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4425|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1001;
  assign _08669_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4424|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 4'b1000;
  assign _08670_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4423|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 3'b111;
  assign _08671_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4422|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 3'b110;
  assign _08672_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4421|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 3'b101;
  assign _08673_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4420|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 3'b100;
  assign _08674_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4419|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 2'b11;
  assign _08675_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4418|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 2'b10;
  assign _08676_ = vec_sum_025_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4417|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4416" *) 1'b1;
  function [7:0] _18170_;
    input [7:0] a;
    input [199:0] b;
    input [24:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *)
    (* parallel_case *)
    casez (s)
      25'b????????????????????????1:
        _18170_ = b[7:0];
      25'b???????????????????????1?:
        _18170_ = b[15:8];
      25'b??????????????????????1??:
        _18170_ = b[23:16];
      25'b?????????????????????1???:
        _18170_ = b[31:24];
      25'b????????????????????1????:
        _18170_ = b[39:32];
      25'b???????????????????1?????:
        _18170_ = b[47:40];
      25'b??????????????????1??????:
        _18170_ = b[55:48];
      25'b?????????????????1???????:
        _18170_ = b[63:56];
      25'b????????????????1????????:
        _18170_ = b[71:64];
      25'b???????????????1?????????:
        _18170_ = b[79:72];
      25'b??????????????1??????????:
        _18170_ = b[87:80];
      25'b?????????????1???????????:
        _18170_ = b[95:88];
      25'b????????????1????????????:
        _18170_ = b[103:96];
      25'b???????????1?????????????:
        _18170_ = b[111:104];
      25'b??????????1??????????????:
        _18170_ = b[119:112];
      25'b?????????1???????????????:
        _18170_ = b[127:120];
      25'b????????1????????????????:
        _18170_ = b[135:128];
      25'b???????1?????????????????:
        _18170_ = b[143:136];
      25'b??????1??????????????????:
        _18170_ = b[151:144];
      25'b?????1???????????????????:
        _18170_ = b[159:152];
      25'b????1????????????????????:
        _18170_ = b[167:160];
      25'b???1?????????????????????:
        _18170_ = b[175:168];
      25'b??1??????????????????????:
        _18170_ = b[183:176];
      25'b?1???????????????????????:
        _18170_ = b[191:184];
      25'b1????????????????????????:
        _18170_ = b[199:192];
      default:
        _18170_ = a;
    endcase
  endfunction
  assign vec_data_024 = _18170_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184], data_d1[199:192] }, { _08701_, _08700_, _08699_, _08698_, _08697_, _08696_, _08695_, _08694_, _08693_, _08692_, _08691_, _08690_, _08689_, _08688_, _08687_, _08686_, _08685_, _08684_, _08683_, _08682_, _08681_, _08680_, _08679_, _08678_, _08677_ });
  assign _08677_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4408|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b11001;
  assign _08678_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4407|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b11000;
  assign _08679_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4406|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10111;
  assign _08680_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4405|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10110;
  assign _08681_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4404|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10101;
  assign _08682_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4403|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10100;
  assign _08683_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4402|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10011;
  assign _08684_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4401|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10010;
  assign _08685_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4400|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10001;
  assign _08686_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4399|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 5'b10000;
  assign _08687_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4398|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1111;
  assign _08688_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4397|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1110;
  assign _08689_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4396|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1101;
  assign _08690_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4395|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1100;
  assign _08691_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4394|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1011;
  assign _08692_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4393|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1010;
  assign _08693_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4392|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1001;
  assign _08694_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4391|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 4'b1000;
  assign _08695_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4390|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 3'b111;
  assign _08696_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4389|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 3'b110;
  assign _08697_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4388|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 3'b101;
  assign _08698_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4387|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 3'b100;
  assign _08699_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4386|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 2'b11;
  assign _08700_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4385|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 2'b10;
  assign _08701_ = vec_sum_024_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4384|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4383" *) 1'b1;
  function [7:0] _18196_;
    input [7:0] a;
    input [191:0] b;
    input [23:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *)
    (* parallel_case *)
    casez (s)
      24'b???????????????????????1:
        _18196_ = b[7:0];
      24'b??????????????????????1?:
        _18196_ = b[15:8];
      24'b?????????????????????1??:
        _18196_ = b[23:16];
      24'b????????????????????1???:
        _18196_ = b[31:24];
      24'b???????????????????1????:
        _18196_ = b[39:32];
      24'b??????????????????1?????:
        _18196_ = b[47:40];
      24'b?????????????????1??????:
        _18196_ = b[55:48];
      24'b????????????????1???????:
        _18196_ = b[63:56];
      24'b???????????????1????????:
        _18196_ = b[71:64];
      24'b??????????????1?????????:
        _18196_ = b[79:72];
      24'b?????????????1??????????:
        _18196_ = b[87:80];
      24'b????????????1???????????:
        _18196_ = b[95:88];
      24'b???????????1????????????:
        _18196_ = b[103:96];
      24'b??????????1?????????????:
        _18196_ = b[111:104];
      24'b?????????1??????????????:
        _18196_ = b[119:112];
      24'b????????1???????????????:
        _18196_ = b[127:120];
      24'b???????1????????????????:
        _18196_ = b[135:128];
      24'b??????1?????????????????:
        _18196_ = b[143:136];
      24'b?????1??????????????????:
        _18196_ = b[151:144];
      24'b????1???????????????????:
        _18196_ = b[159:152];
      24'b???1????????????????????:
        _18196_ = b[167:160];
      24'b??1?????????????????????:
        _18196_ = b[175:168];
      24'b?1??????????????????????:
        _18196_ = b[183:176];
      24'b1???????????????????????:
        _18196_ = b[191:184];
      default:
        _18196_ = a;
    endcase
  endfunction
  assign vec_data_023 = _18196_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176], data_d1[191:184] }, { _08725_, _08724_, _08723_, _08722_, _08721_, _08720_, _08719_, _08718_, _08717_, _08716_, _08715_, _08714_, _08713_, _08712_, _08711_, _08710_, _08709_, _08708_, _08707_, _08706_, _08705_, _08704_, _08703_, _08702_ });
  assign _08702_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4375|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b11000;
  assign _08703_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4374|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10111;
  assign _08704_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4373|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10110;
  assign _08705_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4372|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10101;
  assign _08706_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4371|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10100;
  assign _08707_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4370|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10011;
  assign _08708_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4369|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10010;
  assign _08709_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4368|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10001;
  assign _08710_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4367|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 5'b10000;
  assign _08711_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4366|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1111;
  assign _08712_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4365|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1110;
  assign _08713_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4364|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1101;
  assign _08714_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4363|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1100;
  assign _08715_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4362|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1011;
  assign _08716_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4361|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1010;
  assign _08717_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4360|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1001;
  assign _08718_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4359|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 4'b1000;
  assign _08719_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4358|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 3'b111;
  assign _08720_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4357|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 3'b110;
  assign _08721_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4356|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 3'b101;
  assign _08722_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4355|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 3'b100;
  assign _08723_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4354|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 2'b11;
  assign _08724_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4353|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 2'b10;
  assign _08725_ = vec_sum_023_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4352|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4351" *) 1'b1;
  function [7:0] _18221_;
    input [7:0] a;
    input [183:0] b;
    input [22:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *)
    (* parallel_case *)
    casez (s)
      23'b??????????????????????1:
        _18221_ = b[7:0];
      23'b?????????????????????1?:
        _18221_ = b[15:8];
      23'b????????????????????1??:
        _18221_ = b[23:16];
      23'b???????????????????1???:
        _18221_ = b[31:24];
      23'b??????????????????1????:
        _18221_ = b[39:32];
      23'b?????????????????1?????:
        _18221_ = b[47:40];
      23'b????????????????1??????:
        _18221_ = b[55:48];
      23'b???????????????1???????:
        _18221_ = b[63:56];
      23'b??????????????1????????:
        _18221_ = b[71:64];
      23'b?????????????1?????????:
        _18221_ = b[79:72];
      23'b????????????1??????????:
        _18221_ = b[87:80];
      23'b???????????1???????????:
        _18221_ = b[95:88];
      23'b??????????1????????????:
        _18221_ = b[103:96];
      23'b?????????1?????????????:
        _18221_ = b[111:104];
      23'b????????1??????????????:
        _18221_ = b[119:112];
      23'b???????1???????????????:
        _18221_ = b[127:120];
      23'b??????1????????????????:
        _18221_ = b[135:128];
      23'b?????1?????????????????:
        _18221_ = b[143:136];
      23'b????1??????????????????:
        _18221_ = b[151:144];
      23'b???1???????????????????:
        _18221_ = b[159:152];
      23'b??1????????????????????:
        _18221_ = b[167:160];
      23'b?1?????????????????????:
        _18221_ = b[175:168];
      23'b1??????????????????????:
        _18221_ = b[183:176];
      default:
        _18221_ = a;
    endcase
  endfunction
  assign vec_data_022 = _18221_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168], data_d1[183:176] }, { _08748_, _08747_, _08746_, _08745_, _08744_, _08743_, _08742_, _08741_, _08740_, _08739_, _08738_, _08737_, _08736_, _08735_, _08734_, _08733_, _08732_, _08731_, _08730_, _08729_, _08728_, _08727_, _08726_ });
  assign _08726_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4343|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10111;
  assign _08727_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4342|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10110;
  assign _08728_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4341|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10101;
  assign _08729_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4340|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10100;
  assign _08730_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4339|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10011;
  assign _08731_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4338|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10010;
  assign _08732_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4337|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10001;
  assign _08733_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4336|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 5'b10000;
  assign _08734_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4335|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1111;
  assign _08735_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4334|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1110;
  assign _08736_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4333|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1101;
  assign _08737_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4332|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1100;
  assign _08738_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4331|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1011;
  assign _08739_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4330|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1010;
  assign _08740_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4329|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1001;
  assign _08741_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4328|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 4'b1000;
  assign _08742_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4327|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 3'b111;
  assign _08743_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4326|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 3'b110;
  assign _08744_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4325|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 3'b101;
  assign _08745_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4324|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 3'b100;
  assign _08746_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4323|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 2'b11;
  assign _08747_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4322|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 2'b10;
  assign _08748_ = vec_sum_022_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4321|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4320" *) 1'b1;
  function [7:0] _18245_;
    input [7:0] a;
    input [175:0] b;
    input [21:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *)
    (* parallel_case *)
    casez (s)
      22'b?????????????????????1:
        _18245_ = b[7:0];
      22'b????????????????????1?:
        _18245_ = b[15:8];
      22'b???????????????????1??:
        _18245_ = b[23:16];
      22'b??????????????????1???:
        _18245_ = b[31:24];
      22'b?????????????????1????:
        _18245_ = b[39:32];
      22'b????????????????1?????:
        _18245_ = b[47:40];
      22'b???????????????1??????:
        _18245_ = b[55:48];
      22'b??????????????1???????:
        _18245_ = b[63:56];
      22'b?????????????1????????:
        _18245_ = b[71:64];
      22'b????????????1?????????:
        _18245_ = b[79:72];
      22'b???????????1??????????:
        _18245_ = b[87:80];
      22'b??????????1???????????:
        _18245_ = b[95:88];
      22'b?????????1????????????:
        _18245_ = b[103:96];
      22'b????????1?????????????:
        _18245_ = b[111:104];
      22'b???????1??????????????:
        _18245_ = b[119:112];
      22'b??????1???????????????:
        _18245_ = b[127:120];
      22'b?????1????????????????:
        _18245_ = b[135:128];
      22'b????1?????????????????:
        _18245_ = b[143:136];
      22'b???1??????????????????:
        _18245_ = b[151:144];
      22'b??1???????????????????:
        _18245_ = b[159:152];
      22'b?1????????????????????:
        _18245_ = b[167:160];
      22'b1?????????????????????:
        _18245_ = b[175:168];
      default:
        _18245_ = a;
    endcase
  endfunction
  assign vec_data_021 = _18245_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160], data_d1[175:168] }, { _08770_, _08769_, _08768_, _08767_, _08766_, _08765_, _08764_, _08763_, _08762_, _08761_, _08760_, _08759_, _08758_, _08757_, _08756_, _08755_, _08754_, _08753_, _08752_, _08751_, _08750_, _08749_ });
  assign _08749_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4312|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10110;
  assign _08750_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4311|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10101;
  assign _08751_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4310|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10100;
  assign _08752_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4309|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10011;
  assign _08753_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4308|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10010;
  assign _08754_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4307|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10001;
  assign _08755_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4306|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 5'b10000;
  assign _08756_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4305|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1111;
  assign _08757_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4304|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1110;
  assign _08758_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4303|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1101;
  assign _08759_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4302|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1100;
  assign _08760_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4301|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1011;
  assign _08761_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4300|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1010;
  assign _08762_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4299|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1001;
  assign _08763_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4298|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 4'b1000;
  assign _08764_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4297|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 3'b111;
  assign _08765_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4296|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 3'b110;
  assign _08766_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4295|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 3'b101;
  assign _08767_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4294|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 3'b100;
  assign _08768_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4293|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 2'b11;
  assign _08769_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4292|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 2'b10;
  assign _08770_ = vec_sum_021_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4291|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4290" *) 1'b1;
  function [7:0] _18268_;
    input [7:0] a;
    input [167:0] b;
    input [20:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *)
    (* parallel_case *)
    casez (s)
      21'b????????????????????1:
        _18268_ = b[7:0];
      21'b???????????????????1?:
        _18268_ = b[15:8];
      21'b??????????????????1??:
        _18268_ = b[23:16];
      21'b?????????????????1???:
        _18268_ = b[31:24];
      21'b????????????????1????:
        _18268_ = b[39:32];
      21'b???????????????1?????:
        _18268_ = b[47:40];
      21'b??????????????1??????:
        _18268_ = b[55:48];
      21'b?????????????1???????:
        _18268_ = b[63:56];
      21'b????????????1????????:
        _18268_ = b[71:64];
      21'b???????????1?????????:
        _18268_ = b[79:72];
      21'b??????????1??????????:
        _18268_ = b[87:80];
      21'b?????????1???????????:
        _18268_ = b[95:88];
      21'b????????1????????????:
        _18268_ = b[103:96];
      21'b???????1?????????????:
        _18268_ = b[111:104];
      21'b??????1??????????????:
        _18268_ = b[119:112];
      21'b?????1???????????????:
        _18268_ = b[127:120];
      21'b????1????????????????:
        _18268_ = b[135:128];
      21'b???1?????????????????:
        _18268_ = b[143:136];
      21'b??1??????????????????:
        _18268_ = b[151:144];
      21'b?1???????????????????:
        _18268_ = b[159:152];
      21'b1????????????????????:
        _18268_ = b[167:160];
      default:
        _18268_ = a;
    endcase
  endfunction
  assign vec_data_020 = _18268_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152], data_d1[167:160] }, { _08791_, _08790_, _08789_, _08788_, _08787_, _08786_, _08785_, _08784_, _08783_, _08782_, _08781_, _08780_, _08779_, _08778_, _08777_, _08776_, _08775_, _08774_, _08773_, _08772_, _08771_ });
  assign _08771_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4282|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10101;
  assign _08772_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4281|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10100;
  assign _08773_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4280|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10011;
  assign _08774_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4279|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10010;
  assign _08775_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4278|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10001;
  assign _08776_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4277|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 5'b10000;
  assign _08777_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4276|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1111;
  assign _08778_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4275|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1110;
  assign _08779_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4274|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1101;
  assign _08780_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4273|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1100;
  assign _08781_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4272|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1011;
  assign _08782_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4271|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1010;
  assign _08783_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4270|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1001;
  assign _08784_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4269|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 4'b1000;
  assign _08785_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4268|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 3'b111;
  assign _08786_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4267|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 3'b110;
  assign _08787_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4266|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 3'b101;
  assign _08788_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4265|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 3'b100;
  assign _08789_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4264|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 2'b11;
  assign _08790_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4263|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 2'b10;
  assign _08791_ = vec_sum_020_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4262|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4261" *) 1'b1;
  function [7:0] _18290_;
    input [7:0] a;
    input [159:0] b;
    input [19:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *)
    (* parallel_case *)
    casez (s)
      20'b???????????????????1:
        _18290_ = b[7:0];
      20'b??????????????????1?:
        _18290_ = b[15:8];
      20'b?????????????????1??:
        _18290_ = b[23:16];
      20'b????????????????1???:
        _18290_ = b[31:24];
      20'b???????????????1????:
        _18290_ = b[39:32];
      20'b??????????????1?????:
        _18290_ = b[47:40];
      20'b?????????????1??????:
        _18290_ = b[55:48];
      20'b????????????1???????:
        _18290_ = b[63:56];
      20'b???????????1????????:
        _18290_ = b[71:64];
      20'b??????????1?????????:
        _18290_ = b[79:72];
      20'b?????????1??????????:
        _18290_ = b[87:80];
      20'b????????1???????????:
        _18290_ = b[95:88];
      20'b???????1????????????:
        _18290_ = b[103:96];
      20'b??????1?????????????:
        _18290_ = b[111:104];
      20'b?????1??????????????:
        _18290_ = b[119:112];
      20'b????1???????????????:
        _18290_ = b[127:120];
      20'b???1????????????????:
        _18290_ = b[135:128];
      20'b??1?????????????????:
        _18290_ = b[143:136];
      20'b?1??????????????????:
        _18290_ = b[151:144];
      20'b1???????????????????:
        _18290_ = b[159:152];
      default:
        _18290_ = a;
    endcase
  endfunction
  assign vec_data_019 = _18290_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144], data_d1[159:152] }, { _08811_, _08810_, _08809_, _08808_, _08807_, _08806_, _08805_, _08804_, _08803_, _08802_, _08801_, _08800_, _08799_, _08798_, _08797_, _08796_, _08795_, _08794_, _08793_, _08792_ });
  assign _08792_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4253|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 5'b10100;
  assign _08793_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4252|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 5'b10011;
  assign _08794_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4251|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 5'b10010;
  assign _08795_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4250|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 5'b10001;
  assign _08796_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4249|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 5'b10000;
  assign _08797_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4248|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1111;
  assign _08798_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4247|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1110;
  assign _08799_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4246|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1101;
  assign _08800_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4245|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1100;
  assign _08801_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4244|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1011;
  assign _08802_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4243|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1010;
  assign _08803_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4242|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1001;
  assign _08804_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4241|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 4'b1000;
  assign _08805_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4240|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 3'b111;
  assign _08806_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4239|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 3'b110;
  assign _08807_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4238|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 3'b101;
  assign _08808_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4237|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 3'b100;
  assign _08809_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4236|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 2'b11;
  assign _08810_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4235|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 2'b10;
  assign _08811_ = vec_sum_019_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4234|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4233" *) 1'b1;
  function [7:0] _18311_;
    input [7:0] a;
    input [151:0] b;
    input [18:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *)
    (* parallel_case *)
    casez (s)
      19'b??????????????????1:
        _18311_ = b[7:0];
      19'b?????????????????1?:
        _18311_ = b[15:8];
      19'b????????????????1??:
        _18311_ = b[23:16];
      19'b???????????????1???:
        _18311_ = b[31:24];
      19'b??????????????1????:
        _18311_ = b[39:32];
      19'b?????????????1?????:
        _18311_ = b[47:40];
      19'b????????????1??????:
        _18311_ = b[55:48];
      19'b???????????1???????:
        _18311_ = b[63:56];
      19'b??????????1????????:
        _18311_ = b[71:64];
      19'b?????????1?????????:
        _18311_ = b[79:72];
      19'b????????1??????????:
        _18311_ = b[87:80];
      19'b???????1???????????:
        _18311_ = b[95:88];
      19'b??????1????????????:
        _18311_ = b[103:96];
      19'b?????1?????????????:
        _18311_ = b[111:104];
      19'b????1??????????????:
        _18311_ = b[119:112];
      19'b???1???????????????:
        _18311_ = b[127:120];
      19'b??1????????????????:
        _18311_ = b[135:128];
      19'b?1?????????????????:
        _18311_ = b[143:136];
      19'b1??????????????????:
        _18311_ = b[151:144];
      default:
        _18311_ = a;
    endcase
  endfunction
  assign vec_data_018 = _18311_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136], data_d1[151:144] }, { _08830_, _08829_, _08828_, _08827_, _08826_, _08825_, _08824_, _08823_, _08822_, _08821_, _08820_, _08819_, _08818_, _08817_, _08816_, _08815_, _08814_, _08813_, _08812_ });
  assign _08812_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4225|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 5'b10011;
  assign _08813_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4224|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 5'b10010;
  assign _08814_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4223|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 5'b10001;
  assign _08815_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4222|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 5'b10000;
  assign _08816_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4221|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1111;
  assign _08817_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4220|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1110;
  assign _08818_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4219|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1101;
  assign _08819_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4218|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1100;
  assign _08820_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4217|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1011;
  assign _08821_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4216|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1010;
  assign _08822_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4215|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1001;
  assign _08823_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4214|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 4'b1000;
  assign _08824_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4213|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 3'b111;
  assign _08825_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4212|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 3'b110;
  assign _08826_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4211|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 3'b101;
  assign _08827_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4210|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 3'b100;
  assign _08828_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4209|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 2'b11;
  assign _08829_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4208|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 2'b10;
  assign _08830_ = vec_sum_018_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4207|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4206" *) 1'b1;
  function [7:0] _18331_;
    input [7:0] a;
    input [143:0] b;
    input [17:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *)
    (* parallel_case *)
    casez (s)
      18'b?????????????????1:
        _18331_ = b[7:0];
      18'b????????????????1?:
        _18331_ = b[15:8];
      18'b???????????????1??:
        _18331_ = b[23:16];
      18'b??????????????1???:
        _18331_ = b[31:24];
      18'b?????????????1????:
        _18331_ = b[39:32];
      18'b????????????1?????:
        _18331_ = b[47:40];
      18'b???????????1??????:
        _18331_ = b[55:48];
      18'b??????????1???????:
        _18331_ = b[63:56];
      18'b?????????1????????:
        _18331_ = b[71:64];
      18'b????????1?????????:
        _18331_ = b[79:72];
      18'b???????1??????????:
        _18331_ = b[87:80];
      18'b??????1???????????:
        _18331_ = b[95:88];
      18'b?????1????????????:
        _18331_ = b[103:96];
      18'b????1?????????????:
        _18331_ = b[111:104];
      18'b???1??????????????:
        _18331_ = b[119:112];
      18'b??1???????????????:
        _18331_ = b[127:120];
      18'b?1????????????????:
        _18331_ = b[135:128];
      18'b1?????????????????:
        _18331_ = b[143:136];
      default:
        _18331_ = a;
    endcase
  endfunction
  assign vec_data_017 = _18331_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128], data_d1[143:136] }, { _08848_, _08847_, _08846_, _08845_, _08844_, _08843_, _08842_, _08841_, _08840_, _08839_, _08838_, _08837_, _08836_, _08835_, _08834_, _08833_, _08832_, _08831_ });
  assign _08831_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4198|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 5'b10010;
  assign _08832_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4197|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 5'b10001;
  assign _08833_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4196|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 5'b10000;
  assign _08834_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4195|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1111;
  assign _08835_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4194|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1110;
  assign _08836_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4193|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1101;
  assign _08837_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4192|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1100;
  assign _08838_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4191|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1011;
  assign _08839_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4190|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1010;
  assign _08840_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4189|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1001;
  assign _08841_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4188|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 4'b1000;
  assign _08842_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4187|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 3'b111;
  assign _08843_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4186|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 3'b110;
  assign _08844_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4185|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 3'b101;
  assign _08845_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4184|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 3'b100;
  assign _08846_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4183|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 2'b11;
  assign _08847_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4182|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 2'b10;
  assign _08848_ = vec_sum_017_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4181|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4180" *) 1'b1;
  function [7:0] _18350_;
    input [7:0] a;
    input [135:0] b;
    input [16:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *)
    (* parallel_case *)
    casez (s)
      17'b????????????????1:
        _18350_ = b[7:0];
      17'b???????????????1?:
        _18350_ = b[15:8];
      17'b??????????????1??:
        _18350_ = b[23:16];
      17'b?????????????1???:
        _18350_ = b[31:24];
      17'b????????????1????:
        _18350_ = b[39:32];
      17'b???????????1?????:
        _18350_ = b[47:40];
      17'b??????????1??????:
        _18350_ = b[55:48];
      17'b?????????1???????:
        _18350_ = b[63:56];
      17'b????????1????????:
        _18350_ = b[71:64];
      17'b???????1?????????:
        _18350_ = b[79:72];
      17'b??????1??????????:
        _18350_ = b[87:80];
      17'b?????1???????????:
        _18350_ = b[95:88];
      17'b????1????????????:
        _18350_ = b[103:96];
      17'b???1?????????????:
        _18350_ = b[111:104];
      17'b??1??????????????:
        _18350_ = b[119:112];
      17'b?1???????????????:
        _18350_ = b[127:120];
      17'b1????????????????:
        _18350_ = b[135:128];
      default:
        _18350_ = a;
    endcase
  endfunction
  assign vec_data_016 = _18350_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120], data_d1[135:128] }, { _08865_, _08864_, _08863_, _08862_, _08861_, _08860_, _08859_, _08858_, _08857_, _08856_, _08855_, _08854_, _08853_, _08852_, _08851_, _08850_, _08849_ });
  assign _08849_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4172|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 5'b10001;
  assign _08850_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4171|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 5'b10000;
  assign _08851_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4170|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1111;
  assign _08852_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4169|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1110;
  assign _08853_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4168|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1101;
  assign _08854_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4167|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1100;
  assign _08855_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4166|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1011;
  assign _08856_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4165|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1010;
  assign _08857_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4164|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1001;
  assign _08858_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4163|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 4'b1000;
  assign _08859_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4162|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 3'b111;
  assign _08860_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4161|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 3'b110;
  assign _08861_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4160|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 3'b101;
  assign _08862_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4159|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 3'b100;
  assign _08863_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4158|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 2'b11;
  assign _08864_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4157|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 2'b10;
  assign _08865_ = vec_sum_016_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4156|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4155" *) 1'b1;
  function [7:0] _18368_;
    input [7:0] a;
    input [127:0] b;
    input [15:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *)
    (* parallel_case *)
    casez (s)
      16'b???????????????1:
        _18368_ = b[7:0];
      16'b??????????????1?:
        _18368_ = b[15:8];
      16'b?????????????1??:
        _18368_ = b[23:16];
      16'b????????????1???:
        _18368_ = b[31:24];
      16'b???????????1????:
        _18368_ = b[39:32];
      16'b??????????1?????:
        _18368_ = b[47:40];
      16'b?????????1??????:
        _18368_ = b[55:48];
      16'b????????1???????:
        _18368_ = b[63:56];
      16'b???????1????????:
        _18368_ = b[71:64];
      16'b??????1?????????:
        _18368_ = b[79:72];
      16'b?????1??????????:
        _18368_ = b[87:80];
      16'b????1???????????:
        _18368_ = b[95:88];
      16'b???1????????????:
        _18368_ = b[103:96];
      16'b??1?????????????:
        _18368_ = b[111:104];
      16'b?1??????????????:
        _18368_ = b[119:112];
      16'b1???????????????:
        _18368_ = b[127:120];
      default:
        _18368_ = a;
    endcase
  endfunction
  assign vec_data_015 = _18368_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112], data_d1[127:120] }, { _08881_, _08880_, _08879_, _08878_, _08877_, _08876_, _08875_, _08874_, _08873_, _08872_, _08871_, _08870_, _08869_, _08868_, _08867_, _08866_ });
  assign _08866_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4147|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 5'b10000;
  assign _08867_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4146|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1111;
  assign _08868_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4145|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1110;
  assign _08869_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4144|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1101;
  assign _08870_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4143|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1100;
  assign _08871_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4142|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1011;
  assign _08872_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4141|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1010;
  assign _08873_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4140|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1001;
  assign _08874_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4139|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 4'b1000;
  assign _08875_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4138|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 3'b111;
  assign _08876_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4137|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 3'b110;
  assign _08877_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4136|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 3'b101;
  assign _08878_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4135|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 3'b100;
  assign _08879_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4134|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 2'b11;
  assign _08880_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4133|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 2'b10;
  assign _08881_ = vec_sum_015_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4132|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4131" *) 1'b1;
  function [7:0] _18385_;
    input [7:0] a;
    input [119:0] b;
    input [14:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *)
    (* parallel_case *)
    casez (s)
      15'b??????????????1:
        _18385_ = b[7:0];
      15'b?????????????1?:
        _18385_ = b[15:8];
      15'b????????????1??:
        _18385_ = b[23:16];
      15'b???????????1???:
        _18385_ = b[31:24];
      15'b??????????1????:
        _18385_ = b[39:32];
      15'b?????????1?????:
        _18385_ = b[47:40];
      15'b????????1??????:
        _18385_ = b[55:48];
      15'b???????1???????:
        _18385_ = b[63:56];
      15'b??????1????????:
        _18385_ = b[71:64];
      15'b?????1?????????:
        _18385_ = b[79:72];
      15'b????1??????????:
        _18385_ = b[87:80];
      15'b???1???????????:
        _18385_ = b[95:88];
      15'b??1????????????:
        _18385_ = b[103:96];
      15'b?1?????????????:
        _18385_ = b[111:104];
      15'b1??????????????:
        _18385_ = b[119:112];
      default:
        _18385_ = a;
    endcase
  endfunction
  assign vec_data_014 = _18385_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104], data_d1[119:112] }, { _08896_, _08895_, _08894_, _08893_, _08892_, _08891_, _08890_, _08889_, _08888_, _08887_, _08886_, _08885_, _08884_, _08883_, _08882_ });
  assign _08882_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4123|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1111;
  assign _08883_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4122|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1110;
  assign _08884_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4121|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1101;
  assign _08885_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4120|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1100;
  assign _08886_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4119|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1011;
  assign _08887_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4118|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1010;
  assign _08888_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4117|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1001;
  assign _08889_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4116|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 4'b1000;
  assign _08890_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4115|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 3'b111;
  assign _08891_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4114|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 3'b110;
  assign _08892_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4113|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 3'b101;
  assign _08893_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4112|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 3'b100;
  assign _08894_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4111|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 2'b11;
  assign _08895_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4110|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 2'b10;
  assign _08896_ = vec_sum_014_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4109|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4108" *) 1'b1;
  function [7:0] _18401_;
    input [7:0] a;
    input [111:0] b;
    input [13:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *)
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        _18401_ = b[7:0];
      14'b????????????1?:
        _18401_ = b[15:8];
      14'b???????????1??:
        _18401_ = b[23:16];
      14'b??????????1???:
        _18401_ = b[31:24];
      14'b?????????1????:
        _18401_ = b[39:32];
      14'b????????1?????:
        _18401_ = b[47:40];
      14'b???????1??????:
        _18401_ = b[55:48];
      14'b??????1???????:
        _18401_ = b[63:56];
      14'b?????1????????:
        _18401_ = b[71:64];
      14'b????1?????????:
        _18401_ = b[79:72];
      14'b???1??????????:
        _18401_ = b[87:80];
      14'b??1???????????:
        _18401_ = b[95:88];
      14'b?1????????????:
        _18401_ = b[103:96];
      14'b1?????????????:
        _18401_ = b[111:104];
      default:
        _18401_ = a;
    endcase
  endfunction
  assign vec_data_013 = _18401_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96], data_d1[111:104] }, { _08910_, _08909_, _08908_, _08907_, _08906_, _08905_, _08904_, _08903_, _08902_, _08901_, _08900_, _08899_, _08898_, _08897_ });
  assign _08897_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4100|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1110;
  assign _08898_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4099|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1101;
  assign _08899_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4098|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1100;
  assign _08900_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4097|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1011;
  assign _08901_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4096|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1010;
  assign _08902_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4095|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1001;
  assign _08903_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4094|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 4'b1000;
  assign _08904_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4093|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 3'b111;
  assign _08905_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4092|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 3'b110;
  assign _08906_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4091|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 3'b101;
  assign _08907_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4090|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 3'b100;
  assign _08908_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4089|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 2'b11;
  assign _08909_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4088|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 2'b10;
  assign _08910_ = vec_sum_013_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4087|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4086" *) 1'b1;
  function [7:0] _18416_;
    input [7:0] a;
    input [103:0] b;
    input [12:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *)
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        _18416_ = b[7:0];
      13'b???????????1?:
        _18416_ = b[15:8];
      13'b??????????1??:
        _18416_ = b[23:16];
      13'b?????????1???:
        _18416_ = b[31:24];
      13'b????????1????:
        _18416_ = b[39:32];
      13'b???????1?????:
        _18416_ = b[47:40];
      13'b??????1??????:
        _18416_ = b[55:48];
      13'b?????1???????:
        _18416_ = b[63:56];
      13'b????1????????:
        _18416_ = b[71:64];
      13'b???1?????????:
        _18416_ = b[79:72];
      13'b??1??????????:
        _18416_ = b[87:80];
      13'b?1???????????:
        _18416_ = b[95:88];
      13'b1????????????:
        _18416_ = b[103:96];
      default:
        _18416_ = a;
    endcase
  endfunction
  assign vec_data_012 = _18416_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88], data_d1[103:96] }, { _08923_, _08922_, _08921_, _08920_, _08919_, _08918_, _08917_, _08916_, _08915_, _08914_, _08913_, _08912_, _08911_ });
  assign _08911_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4078|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1101;
  assign _08912_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4077|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1100;
  assign _08913_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4076|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1011;
  assign _08914_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4075|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1010;
  assign _08915_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4074|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1001;
  assign _08916_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4073|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 4'b1000;
  assign _08917_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4072|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 3'b111;
  assign _08918_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4071|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 3'b110;
  assign _08919_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4070|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 3'b101;
  assign _08920_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4069|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 3'b100;
  assign _08921_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4068|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 2'b11;
  assign _08922_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4067|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 2'b10;
  assign _08923_ = vec_sum_012_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4066|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4065" *) 1'b1;
  function [7:0] _18430_;
    input [7:0] a;
    input [95:0] b;
    input [11:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *)
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        _18430_ = b[7:0];
      12'b??????????1?:
        _18430_ = b[15:8];
      12'b?????????1??:
        _18430_ = b[23:16];
      12'b????????1???:
        _18430_ = b[31:24];
      12'b???????1????:
        _18430_ = b[39:32];
      12'b??????1?????:
        _18430_ = b[47:40];
      12'b?????1??????:
        _18430_ = b[55:48];
      12'b????1???????:
        _18430_ = b[63:56];
      12'b???1????????:
        _18430_ = b[71:64];
      12'b??1?????????:
        _18430_ = b[79:72];
      12'b?1??????????:
        _18430_ = b[87:80];
      12'b1???????????:
        _18430_ = b[95:88];
      default:
        _18430_ = a;
    endcase
  endfunction
  assign vec_data_011 = _18430_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80], data_d1[95:88] }, { _08935_, _08934_, _08933_, _08932_, _08931_, _08930_, _08929_, _08928_, _08927_, _08926_, _08925_, _08924_ });
  assign _08924_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4057|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 4'b1100;
  assign _08925_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4056|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 4'b1011;
  assign _08926_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4055|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 4'b1010;
  assign _08927_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4054|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 4'b1001;
  assign _08928_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4053|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 4'b1000;
  assign _08929_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4052|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 3'b111;
  assign _08930_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4051|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 3'b110;
  assign _08931_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4050|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 3'b101;
  assign _08932_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4049|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 3'b100;
  assign _08933_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4048|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 2'b11;
  assign _08934_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4047|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 2'b10;
  assign _08935_ = vec_sum_011_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4046|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4045" *) 1'b1;
  function [7:0] _18443_;
    input [7:0] a;
    input [87:0] b;
    input [10:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *)
    (* parallel_case *)
    casez (s)
      11'b??????????1:
        _18443_ = b[7:0];
      11'b?????????1?:
        _18443_ = b[15:8];
      11'b????????1??:
        _18443_ = b[23:16];
      11'b???????1???:
        _18443_ = b[31:24];
      11'b??????1????:
        _18443_ = b[39:32];
      11'b?????1?????:
        _18443_ = b[47:40];
      11'b????1??????:
        _18443_ = b[55:48];
      11'b???1???????:
        _18443_ = b[63:56];
      11'b??1????????:
        _18443_ = b[71:64];
      11'b?1?????????:
        _18443_ = b[79:72];
      11'b1??????????:
        _18443_ = b[87:80];
      default:
        _18443_ = a;
    endcase
  endfunction
  assign vec_data_010 = _18443_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72], data_d1[87:80] }, { _08946_, _08945_, _08944_, _08943_, _08942_, _08941_, _08940_, _08939_, _08938_, _08937_, _08936_ });
  assign _08936_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4037|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 4'b1011;
  assign _08937_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4036|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 4'b1010;
  assign _08938_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4035|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 4'b1001;
  assign _08939_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4034|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 4'b1000;
  assign _08940_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4033|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 3'b111;
  assign _08941_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4032|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 3'b110;
  assign _08942_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4031|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 3'b101;
  assign _08943_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4030|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 3'b100;
  assign _08944_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4029|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 2'b11;
  assign _08945_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4028|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 2'b10;
  assign _08946_ = vec_sum_010_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4027|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4026" *) 1'b1;
  function [7:0] _18455_;
    input [7:0] a;
    input [79:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _18455_ = b[7:0];
      10'b????????1?:
        _18455_ = b[15:8];
      10'b???????1??:
        _18455_ = b[23:16];
      10'b??????1???:
        _18455_ = b[31:24];
      10'b?????1????:
        _18455_ = b[39:32];
      10'b????1?????:
        _18455_ = b[47:40];
      10'b???1??????:
        _18455_ = b[55:48];
      10'b??1???????:
        _18455_ = b[63:56];
      10'b?1????????:
        _18455_ = b[71:64];
      10'b1?????????:
        _18455_ = b[79:72];
      default:
        _18455_ = a;
    endcase
  endfunction
  assign vec_data_009 = _18455_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64], data_d1[79:72] }, { _08956_, _08955_, _08954_, _08953_, _08952_, _08951_, _08950_, _08949_, _08948_, _08947_ });
  assign _08947_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4018|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 4'b1010;
  assign _08948_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4017|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 4'b1001;
  assign _08949_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4016|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 4'b1000;
  assign _08950_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4015|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 3'b111;
  assign _08951_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4014|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 3'b110;
  assign _08952_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4013|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 3'b101;
  assign _08953_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4012|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 3'b100;
  assign _08954_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4011|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 2'b11;
  assign _08955_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4010|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 2'b10;
  assign _08956_ = vec_sum_009_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4009|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4008" *) 1'b1;
  function [7:0] _18466_;
    input [7:0] a;
    input [71:0] b;
    input [8:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *)
    (* parallel_case *)
    casez (s)
      9'b????????1:
        _18466_ = b[7:0];
      9'b???????1?:
        _18466_ = b[15:8];
      9'b??????1??:
        _18466_ = b[23:16];
      9'b?????1???:
        _18466_ = b[31:24];
      9'b????1????:
        _18466_ = b[39:32];
      9'b???1?????:
        _18466_ = b[47:40];
      9'b??1??????:
        _18466_ = b[55:48];
      9'b?1???????:
        _18466_ = b[63:56];
      9'b1????????:
        _18466_ = b[71:64];
      default:
        _18466_ = a;
    endcase
  endfunction
  assign vec_data_008 = _18466_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56], data_d1[71:64] }, { _08965_, _08964_, _08963_, _08962_, _08961_, _08960_, _08959_, _08958_, _08957_ });
  assign _08957_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:4000|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 4'b1001;
  assign _08958_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3999|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 4'b1000;
  assign _08959_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3998|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 3'b111;
  assign _08960_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3997|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 3'b110;
  assign _08961_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3996|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 3'b101;
  assign _08962_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3995|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 3'b100;
  assign _08963_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3994|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 2'b11;
  assign _08964_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3993|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 2'b10;
  assign _08965_ = vec_sum_008_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3992|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3991" *) 1'b1;
  function [7:0] _18476_;
    input [7:0] a;
    input [63:0] b;
    input [7:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *)
    (* parallel_case *)
    casez (s)
      8'b???????1:
        _18476_ = b[7:0];
      8'b??????1?:
        _18476_ = b[15:8];
      8'b?????1??:
        _18476_ = b[23:16];
      8'b????1???:
        _18476_ = b[31:24];
      8'b???1????:
        _18476_ = b[39:32];
      8'b??1?????:
        _18476_ = b[47:40];
      8'b?1??????:
        _18476_ = b[55:48];
      8'b1???????:
        _18476_ = b[63:56];
      default:
        _18476_ = a;
    endcase
  endfunction
  assign vec_data_007 = _18476_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48], data_d1[63:56] }, { _08973_, _08972_, _08971_, _08970_, _08969_, _08968_, _08967_, _08966_ });
  assign _08966_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3983|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 4'b1000;
  assign _08967_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3982|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 3'b111;
  assign _08968_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3981|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 3'b110;
  assign _08969_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3980|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 3'b101;
  assign _08970_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3979|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 3'b100;
  assign _08971_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3978|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 2'b11;
  assign _08972_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3977|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 2'b10;
  assign _08973_ = vec_sum_007_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3976|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3975" *) 1'b1;
  function [7:0] _18485_;
    input [7:0] a;
    input [55:0] b;
    input [6:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *)
    (* parallel_case *)
    casez (s)
      7'b??????1:
        _18485_ = b[7:0];
      7'b?????1?:
        _18485_ = b[15:8];
      7'b????1??:
        _18485_ = b[23:16];
      7'b???1???:
        _18485_ = b[31:24];
      7'b??1????:
        _18485_ = b[39:32];
      7'b?1?????:
        _18485_ = b[47:40];
      7'b1??????:
        _18485_ = b[55:48];
      default:
        _18485_ = a;
    endcase
  endfunction
  assign vec_data_006 = _18485_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40], data_d1[55:48] }, { _08980_, _08979_, _08978_, _08977_, _08976_, _08975_, _08974_ });
  assign _08974_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3967|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 3'b111;
  assign _08975_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3966|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 3'b110;
  assign _08976_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3965|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 3'b101;
  assign _08977_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3964|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 3'b100;
  assign _08978_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3963|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 2'b11;
  assign _08979_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3962|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 2'b10;
  assign _08980_ = vec_sum_006_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3961|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3960" *) 1'b1;
  function [7:0] _18493_;
    input [7:0] a;
    input [47:0] b;
    input [5:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *)
    (* parallel_case *)
    casez (s)
      6'b?????1:
        _18493_ = b[7:0];
      6'b????1?:
        _18493_ = b[15:8];
      6'b???1??:
        _18493_ = b[23:16];
      6'b??1???:
        _18493_ = b[31:24];
      6'b?1????:
        _18493_ = b[39:32];
      6'b1?????:
        _18493_ = b[47:40];
      default:
        _18493_ = a;
    endcase
  endfunction
  assign vec_data_005 = _18493_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32], data_d1[47:40] }, { _08986_, _08985_, _08984_, _08983_, _08982_, _08981_ });
  assign _08981_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3952|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 3'b110;
  assign _08982_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3951|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 3'b101;
  assign _08983_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3950|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 3'b100;
  assign _08984_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3949|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 2'b11;
  assign _08985_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3948|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 2'b10;
  assign _08986_ = vec_sum_005_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3947|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3946" *) 1'b1;
  function [7:0] _18500_;
    input [7:0] a;
    input [39:0] b;
    input [4:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *)
    (* parallel_case *)
    casez (s)
      5'b????1:
        _18500_ = b[7:0];
      5'b???1?:
        _18500_ = b[15:8];
      5'b??1??:
        _18500_ = b[23:16];
      5'b?1???:
        _18500_ = b[31:24];
      5'b1????:
        _18500_ = b[39:32];
      default:
        _18500_ = a;
    endcase
  endfunction
  assign vec_data_004 = _18500_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24], data_d1[39:32] }, { _08991_, _08990_, _08989_, _08988_, _08987_ });
  assign _08987_ = vec_sum_004_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3938|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *) 3'b101;
  assign _08988_ = vec_sum_004_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3937|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *) 3'b100;
  assign _08989_ = vec_sum_004_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3936|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *) 2'b11;
  assign _08990_ = vec_sum_004_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3935|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *) 2'b10;
  assign _08991_ = vec_sum_004_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3934|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3933" *) 1'b1;
  function [7:0] _18506_;
    input [7:0] a;
    input [31:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3921" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _18506_ = b[7:0];
      4'b??1?:
        _18506_ = b[15:8];
      4'b?1??:
        _18506_ = b[23:16];
      4'b1???:
        _18506_ = b[31:24];
      default:
        _18506_ = a;
    endcase
  endfunction
  assign vec_data_003 = _18506_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16], data_d1[31:24] }, { _08995_, _08994_, _08993_, _08992_ });
  assign _08992_ = vec_sum_003_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3925|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3921" *) 3'b100;
  assign _08993_ = vec_sum_003_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3924|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3921" *) 2'b11;
  assign _08994_ = vec_sum_003_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3923|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3921" *) 2'b10;
  assign _08995_ = vec_sum_003_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3922|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3921" *) 1'b1;
  function [7:0] _18511_;
    input [7:0] a;
    input [23:0] b;
    input [2:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3910" *)
    (* parallel_case *)
    casez (s)
      3'b??1:
        _18511_ = b[7:0];
      3'b?1?:
        _18511_ = b[15:8];
      3'b1??:
        _18511_ = b[23:16];
      default:
        _18511_ = a;
    endcase
  endfunction
  assign vec_data_002 = _18511_(8'b00000000, { data_d1[7:0], data_d1[15:8], data_d1[23:16] }, { _08998_, _08997_, _08996_ });
  assign _08996_ = vec_sum_002_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3913|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3910" *) 2'b11;
  assign _08997_ = vec_sum_002_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3912|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3910" *) 2'b10;
  assign _08998_ = vec_sum_002_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3911|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3910" *) 1'b1;
  function [7:0] _18515_;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3900" *)
    (* parallel_case *)
    casez (s)
      2'b?1:
        _18515_ = b[7:0];
      2'b1?:
        _18515_ = b[15:8];
      default:
        _18515_ = a;
    endcase
  endfunction
  assign vec_data_001 = _18515_(8'b00000000, { data_d1[7:0], data_d1[15:8] }, { _09000_, _08999_ });
  assign _08999_ = vec_sum_001_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3902|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3900" *) 2'b10;
  assign _09000_ = vec_sum_001_d1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3901|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3900" *) 1'b1;
  assign vec_data_000 = vec_sum_000_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3892|./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3891" *) data_d1[7:0] : 8'b00000000;
  assign _00389_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3876" *) vec_sum_127 : { _00745_[7], vec_sum_127_d1 };
  assign _00388_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3866" *) vec_sum_126 : vec_sum_126_d1;
  assign _00387_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3856" *) vec_sum_125 : vec_sum_125_d1;
  assign _00386_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3846" *) vec_sum_124 : vec_sum_124_d1;
  assign _00385_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3836" *) vec_sum_123 : vec_sum_123_d1;
  assign _00384_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3826" *) vec_sum_122 : vec_sum_122_d1;
  assign _00383_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3816" *) vec_sum_121 : vec_sum_121_d1;
  assign _00382_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3806" *) vec_sum_120 : vec_sum_120_d1;
  assign _00381_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3796" *) vec_sum_119 : vec_sum_119_d1;
  assign _00380_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3786" *) vec_sum_118 : vec_sum_118_d1;
  assign _00379_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3776" *) vec_sum_117 : vec_sum_117_d1;
  assign _00378_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3766" *) vec_sum_116 : vec_sum_116_d1;
  assign _00377_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3756" *) vec_sum_115 : vec_sum_115_d1;
  assign _00376_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3746" *) vec_sum_114 : vec_sum_114_d1;
  assign _00375_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3736" *) vec_sum_113 : vec_sum_113_d1;
  assign _00374_ = _00744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3726" *) vec_sum_112 : vec_sum_112_d1;
  assign _00373_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3716" *) vec_sum_111 : vec_sum_111_d1;
  assign _00372_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3706" *) vec_sum_110 : vec_sum_110_d1;
  assign _00371_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3696" *) vec_sum_109 : vec_sum_109_d1;
  assign _00370_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3686" *) vec_sum_108 : vec_sum_108_d1;
  assign _00369_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3676" *) vec_sum_107 : vec_sum_107_d1;
  assign _00368_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3666" *) vec_sum_106 : vec_sum_106_d1;
  assign _00367_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3656" *) vec_sum_105 : vec_sum_105_d1;
  assign _00366_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3646" *) vec_sum_104 : vec_sum_104_d1;
  assign _00365_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3636" *) vec_sum_103 : vec_sum_103_d1;
  assign _00364_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3626" *) vec_sum_102 : vec_sum_102_d1;
  assign _00363_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3616" *) vec_sum_101 : vec_sum_101_d1;
  assign _00362_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3606" *) vec_sum_100 : vec_sum_100_d1;
  assign _00361_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3596" *) vec_sum_099 : vec_sum_099_d1;
  assign _00360_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3586" *) vec_sum_098 : vec_sum_098_d1;
  assign _00359_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3576" *) vec_sum_097 : vec_sum_097_d1;
  assign _00358_ = _00743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3566" *) vec_sum_096 : vec_sum_096_d1;
  assign _00357_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3556" *) vec_sum_095 : vec_sum_095_d1;
  assign _00356_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3546" *) vec_sum_094 : vec_sum_094_d1;
  assign _00355_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3536" *) vec_sum_093 : vec_sum_093_d1;
  assign _00354_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3526" *) vec_sum_092 : vec_sum_092_d1;
  assign _00353_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3516" *) vec_sum_091 : vec_sum_091_d1;
  assign _00352_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3506" *) vec_sum_090 : vec_sum_090_d1;
  assign _00351_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3496" *) vec_sum_089 : vec_sum_089_d1;
  assign _00350_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3486" *) vec_sum_088 : vec_sum_088_d1;
  assign _00349_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3476" *) vec_sum_087 : vec_sum_087_d1;
  assign _00348_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3466" *) vec_sum_086 : vec_sum_086_d1;
  assign _00347_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3456" *) vec_sum_085 : vec_sum_085_d1;
  assign _00346_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3446" *) vec_sum_084 : vec_sum_084_d1;
  assign _00345_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3436" *) vec_sum_083 : vec_sum_083_d1;
  assign _00344_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3426" *) vec_sum_082 : vec_sum_082_d1;
  assign _00343_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3416" *) vec_sum_081 : vec_sum_081_d1;
  assign _00342_ = _00742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3406" *) vec_sum_080 : vec_sum_080_d1;
  assign _00341_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3396" *) vec_sum_079 : vec_sum_079_d1;
  assign _00340_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3386" *) vec_sum_078 : vec_sum_078_d1;
  assign _00339_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3376" *) vec_sum_077 : vec_sum_077_d1;
  assign _00338_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3366" *) vec_sum_076 : vec_sum_076_d1;
  assign _00337_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3356" *) vec_sum_075 : vec_sum_075_d1;
  assign _00336_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3346" *) vec_sum_074 : vec_sum_074_d1;
  assign _00335_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3336" *) vec_sum_073 : vec_sum_073_d1;
  assign _00334_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3326" *) vec_sum_072 : vec_sum_072_d1;
  assign _00333_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3316" *) vec_sum_071 : vec_sum_071_d1;
  assign _00332_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3306" *) vec_sum_070 : vec_sum_070_d1;
  assign _00331_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3296" *) vec_sum_069 : vec_sum_069_d1;
  assign _00330_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3286" *) vec_sum_068 : vec_sum_068_d1;
  assign _00329_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3276" *) vec_sum_067 : vec_sum_067_d1;
  assign _00328_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3266" *) vec_sum_066 : vec_sum_066_d1;
  assign _00327_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3256" *) vec_sum_065 : vec_sum_065_d1;
  assign _00326_ = _00741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3246" *) vec_sum_064 : vec_sum_064_d1;
  assign _00325_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3236" *) vec_sum_063 : vec_sum_063_d1;
  assign _00324_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3226" *) vec_sum_062 : vec_sum_062_d1;
  assign _00323_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3216" *) vec_sum_061 : vec_sum_061_d1;
  assign _00322_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3206" *) vec_sum_060 : vec_sum_060_d1;
  assign _00321_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3196" *) vec_sum_059 : vec_sum_059_d1;
  assign _00320_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3186" *) vec_sum_058 : vec_sum_058_d1;
  assign _00319_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3176" *) vec_sum_057 : vec_sum_057_d1;
  assign _00318_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3166" *) vec_sum_056 : vec_sum_056_d1;
  assign _00317_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3156" *) vec_sum_055 : vec_sum_055_d1;
  assign _00316_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3146" *) vec_sum_054 : vec_sum_054_d1;
  assign _00315_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3136" *) vec_sum_053 : vec_sum_053_d1;
  assign _00314_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3126" *) vec_sum_052 : vec_sum_052_d1;
  assign _00313_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3116" *) vec_sum_051 : vec_sum_051_d1;
  assign _00312_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3106" *) vec_sum_050 : vec_sum_050_d1;
  assign _00311_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3096" *) vec_sum_049 : vec_sum_049_d1;
  assign _00310_ = _00740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3086" *) vec_sum_048 : vec_sum_048_d1;
  assign _00309_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3076" *) vec_sum_047 : vec_sum_047_d1;
  assign _00308_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3066" *) vec_sum_046 : vec_sum_046_d1;
  assign _00307_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3056" *) vec_sum_045 : vec_sum_045_d1;
  assign _00306_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3046" *) vec_sum_044 : vec_sum_044_d1;
  assign _00305_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3036" *) vec_sum_043 : vec_sum_043_d1;
  assign _00304_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3026" *) vec_sum_042 : vec_sum_042_d1;
  assign _00303_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3016" *) vec_sum_041 : vec_sum_041_d1;
  assign _00302_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:3006" *) vec_sum_040 : vec_sum_040_d1;
  assign _00301_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2996" *) vec_sum_039 : vec_sum_039_d1;
  assign _00300_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2986" *) vec_sum_038 : vec_sum_038_d1;
  assign _00299_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2976" *) vec_sum_037 : vec_sum_037_d1;
  assign _00298_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2966" *) vec_sum_036 : vec_sum_036_d1;
  assign _00297_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2956" *) vec_sum_035 : vec_sum_035_d1;
  assign _00296_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2946" *) vec_sum_034 : vec_sum_034_d1;
  assign _00295_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2936" *) vec_sum_033 : vec_sum_033_d1;
  assign _00294_ = _00739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2926" *) vec_sum_032 : vec_sum_032_d1;
  assign _00293_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2916" *) vec_sum_031 : vec_sum_031_d1;
  assign _00292_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2906" *) vec_sum_030 : vec_sum_030_d1;
  assign _00291_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2896" *) vec_sum_029 : vec_sum_029_d1;
  assign _00290_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2886" *) vec_sum_028 : vec_sum_028_d1;
  assign _00289_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2876" *) vec_sum_027 : vec_sum_027_d1;
  assign _00288_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2866" *) vec_sum_026 : vec_sum_026_d1;
  assign _00287_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2856" *) vec_sum_025 : vec_sum_025_d1;
  assign _00286_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2846" *) vec_sum_024 : vec_sum_024_d1;
  assign _00285_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2836" *) vec_sum_023 : vec_sum_023_d1;
  assign _00284_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2826" *) vec_sum_022 : vec_sum_022_d1;
  assign _00283_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2816" *) vec_sum_021 : vec_sum_021_d1;
  assign _00282_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2806" *) vec_sum_020 : vec_sum_020_d1;
  assign _00281_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2796" *) vec_sum_019 : vec_sum_019_d1;
  assign _00280_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2786" *) vec_sum_018 : vec_sum_018_d1;
  assign _00279_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2776" *) vec_sum_017 : vec_sum_017_d1;
  assign _00278_ = _00738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2766" *) vec_sum_016 : vec_sum_016_d1;
  assign _00277_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2756" *) vec_sum_015 : vec_sum_015_d1;
  assign _00276_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2746" *) vec_sum_014 : vec_sum_014_d1;
  assign _00275_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2736" *) vec_sum_013 : vec_sum_013_d1;
  assign _00274_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2726" *) vec_sum_012 : vec_sum_012_d1;
  assign _00273_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2716" *) vec_sum_011 : vec_sum_011_d1;
  assign _00272_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2706" *) vec_sum_010 : vec_sum_010_d1;
  assign _00271_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2696" *) vec_sum_009 : vec_sum_009_d1;
  assign _00270_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2686" *) vec_sum_008 : vec_sum_008_d1;
  assign _00269_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2676" *) vec_sum_007 : vec_sum_007_d1;
  assign _00268_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2666" *) vec_sum_006 : vec_sum_006_d1;
  assign _00267_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2656" *) vec_sum_005 : vec_sum_005_d1;
  assign _00266_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2646" *) vec_sum_004 : vec_sum_004_d1;
  assign _00265_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2636" *) vec_sum_003 : vec_sum_003_d1;
  assign _00264_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2626" *) vec_sum_002 : vec_sum_002_d1;
  assign _00263_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2616" *) vec_sum_001 : vec_sum_001_d1;
  assign _00262_ = _00737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2606" *) input_mask_gated[0] : vec_sum_000_d1;
  assign _00003_ = input_pipe_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2596" *) input_sel : sel_d1;
  assign _00001_ = input_mask_en[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2586" *) input_mask : mask_d1;
  assign _00000_ = input_pipe_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:2576" *) input_data : data_d1;
  assign mask_d2_int8_w[0] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20611" *) { vec_data_000_d2[0], vec_data_000_d2[1], vec_data_000_d2[2], vec_data_000_d2[3], vec_data_000_d2[4], vec_data_000_d2[5], vec_data_000_d2[6], vec_data_000_d2[7] };
  assign mask_d2_int8_w[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20612" *) { vec_data_001_d2[0], vec_data_001_d2[1], vec_data_001_d2[2], vec_data_001_d2[3], vec_data_001_d2[4], vec_data_001_d2[5], vec_data_001_d2[6], vec_data_001_d2[7] };
  assign mask_d2_int8_w[2] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20613" *) { vec_data_002_d2[0], vec_data_002_d2[1], vec_data_002_d2[2], vec_data_002_d2[3], vec_data_002_d2[4], vec_data_002_d2[5], vec_data_002_d2[6], vec_data_002_d2[7] };
  assign mask_d2_int8_w[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20614" *) { vec_data_003_d2[0], vec_data_003_d2[1], vec_data_003_d2[2], vec_data_003_d2[3], vec_data_003_d2[4], vec_data_003_d2[5], vec_data_003_d2[6], vec_data_003_d2[7] };
  assign mask_d2_int8_w[4] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20615" *) { vec_data_004_d2[0], vec_data_004_d2[1], vec_data_004_d2[2], vec_data_004_d2[3], vec_data_004_d2[4], vec_data_004_d2[5], vec_data_004_d2[6], vec_data_004_d2[7] };
  assign mask_d2_int8_w[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20616" *) { vec_data_005_d2[0], vec_data_005_d2[1], vec_data_005_d2[2], vec_data_005_d2[3], vec_data_005_d2[4], vec_data_005_d2[5], vec_data_005_d2[6], vec_data_005_d2[7] };
  assign mask_d2_int8_w[6] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20617" *) { vec_data_006_d2[0], vec_data_006_d2[1], vec_data_006_d2[2], vec_data_006_d2[3], vec_data_006_d2[4], vec_data_006_d2[5], vec_data_006_d2[6], vec_data_006_d2[7] };
  assign mask_d2_int8_w[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20618" *) { vec_data_007_d2[0], vec_data_007_d2[1], vec_data_007_d2[2], vec_data_007_d2[3], vec_data_007_d2[4], vec_data_007_d2[5], vec_data_007_d2[6], vec_data_007_d2[7] };
  assign mask_d2_int8_w[8] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20619" *) { vec_data_008_d2[0], vec_data_008_d2[1], vec_data_008_d2[2], vec_data_008_d2[3], vec_data_008_d2[4], vec_data_008_d2[5], vec_data_008_d2[6], vec_data_008_d2[7] };
  assign mask_d2_int8_w[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20620" *) { vec_data_009_d2[0], vec_data_009_d2[1], vec_data_009_d2[2], vec_data_009_d2[3], vec_data_009_d2[4], vec_data_009_d2[5], vec_data_009_d2[6], vec_data_009_d2[7] };
  assign mask_d2_int8_w[10] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20621" *) { vec_data_010_d2[0], vec_data_010_d2[1], vec_data_010_d2[2], vec_data_010_d2[3], vec_data_010_d2[4], vec_data_010_d2[5], vec_data_010_d2[6], vec_data_010_d2[7] };
  assign mask_d2_int8_w[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20622" *) { vec_data_011_d2[0], vec_data_011_d2[1], vec_data_011_d2[2], vec_data_011_d2[3], vec_data_011_d2[4], vec_data_011_d2[5], vec_data_011_d2[6], vec_data_011_d2[7] };
  assign mask_d2_int8_w[12] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20623" *) { vec_data_012_d2[0], vec_data_012_d2[1], vec_data_012_d2[2], vec_data_012_d2[3], vec_data_012_d2[4], vec_data_012_d2[5], vec_data_012_d2[6], vec_data_012_d2[7] };
  assign mask_d2_int8_w[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20624" *) { vec_data_013_d2[0], vec_data_013_d2[1], vec_data_013_d2[2], vec_data_013_d2[3], vec_data_013_d2[4], vec_data_013_d2[5], vec_data_013_d2[6], vec_data_013_d2[7] };
  assign mask_d2_int8_w[14] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20625" *) { vec_data_014_d2[0], vec_data_014_d2[1], vec_data_014_d2[2], vec_data_014_d2[3], vec_data_014_d2[4], vec_data_014_d2[5], vec_data_014_d2[6], vec_data_014_d2[7] };
  assign mask_d2_int8_w[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20626" *) { vec_data_015_d2[0], vec_data_015_d2[1], vec_data_015_d2[2], vec_data_015_d2[3], vec_data_015_d2[4], vec_data_015_d2[5], vec_data_015_d2[6], vec_data_015_d2[7] };
  assign mask_d2_int8_w[16] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20627" *) { vec_data_016_d2[0], vec_data_016_d2[1], vec_data_016_d2[2], vec_data_016_d2[3], vec_data_016_d2[4], vec_data_016_d2[5], vec_data_016_d2[6], vec_data_016_d2[7] };
  assign mask_d2_int8_w[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20628" *) { vec_data_017_d2[0], vec_data_017_d2[1], vec_data_017_d2[2], vec_data_017_d2[3], vec_data_017_d2[4], vec_data_017_d2[5], vec_data_017_d2[6], vec_data_017_d2[7] };
  assign mask_d2_int8_w[18] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20629" *) { vec_data_018_d2[0], vec_data_018_d2[1], vec_data_018_d2[2], vec_data_018_d2[3], vec_data_018_d2[4], vec_data_018_d2[5], vec_data_018_d2[6], vec_data_018_d2[7] };
  assign mask_d2_int8_w[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20630" *) { vec_data_019_d2[0], vec_data_019_d2[1], vec_data_019_d2[2], vec_data_019_d2[3], vec_data_019_d2[4], vec_data_019_d2[5], vec_data_019_d2[6], vec_data_019_d2[7] };
  assign mask_d2_int8_w[20] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20631" *) { vec_data_020_d2[0], vec_data_020_d2[1], vec_data_020_d2[2], vec_data_020_d2[3], vec_data_020_d2[4], vec_data_020_d2[5], vec_data_020_d2[6], vec_data_020_d2[7] };
  assign mask_d2_int8_w[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20632" *) { vec_data_021_d2[0], vec_data_021_d2[1], vec_data_021_d2[2], vec_data_021_d2[3], vec_data_021_d2[4], vec_data_021_d2[5], vec_data_021_d2[6], vec_data_021_d2[7] };
  assign mask_d2_int8_w[22] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20633" *) { vec_data_022_d2[0], vec_data_022_d2[1], vec_data_022_d2[2], vec_data_022_d2[3], vec_data_022_d2[4], vec_data_022_d2[5], vec_data_022_d2[6], vec_data_022_d2[7] };
  assign mask_d2_int8_w[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20634" *) { vec_data_023_d2[0], vec_data_023_d2[1], vec_data_023_d2[2], vec_data_023_d2[3], vec_data_023_d2[4], vec_data_023_d2[5], vec_data_023_d2[6], vec_data_023_d2[7] };
  assign mask_d2_int8_w[24] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20635" *) { vec_data_024_d2[0], vec_data_024_d2[1], vec_data_024_d2[2], vec_data_024_d2[3], vec_data_024_d2[4], vec_data_024_d2[5], vec_data_024_d2[6], vec_data_024_d2[7] };
  assign mask_d2_int8_w[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20636" *) { vec_data_025_d2[0], vec_data_025_d2[1], vec_data_025_d2[2], vec_data_025_d2[3], vec_data_025_d2[4], vec_data_025_d2[5], vec_data_025_d2[6], vec_data_025_d2[7] };
  assign mask_d2_int8_w[26] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20637" *) { vec_data_026_d2[0], vec_data_026_d2[1], vec_data_026_d2[2], vec_data_026_d2[3], vec_data_026_d2[4], vec_data_026_d2[5], vec_data_026_d2[6], vec_data_026_d2[7] };
  assign mask_d2_int8_w[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20638" *) { vec_data_027_d2[0], vec_data_027_d2[1], vec_data_027_d2[2], vec_data_027_d2[3], vec_data_027_d2[4], vec_data_027_d2[5], vec_data_027_d2[6], vec_data_027_d2[7] };
  assign mask_d2_int8_w[28] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20639" *) { vec_data_028_d2[0], vec_data_028_d2[1], vec_data_028_d2[2], vec_data_028_d2[3], vec_data_028_d2[4], vec_data_028_d2[5], vec_data_028_d2[6], vec_data_028_d2[7] };
  assign mask_d2_int8_w[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20640" *) { vec_data_029_d2[0], vec_data_029_d2[1], vec_data_029_d2[2], vec_data_029_d2[3], vec_data_029_d2[4], vec_data_029_d2[5], vec_data_029_d2[6], vec_data_029_d2[7] };
  assign mask_d2_int8_w[30] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20641" *) { vec_data_030_d2[0], vec_data_030_d2[1], vec_data_030_d2[2], vec_data_030_d2[3], vec_data_030_d2[4], vec_data_030_d2[5], vec_data_030_d2[6], vec_data_030_d2[7] };
  assign mask_d2_int8_w[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20642" *) { vec_data_031_d2[0], vec_data_031_d2[1], vec_data_031_d2[2], vec_data_031_d2[3], vec_data_031_d2[4], vec_data_031_d2[5], vec_data_031_d2[6], vec_data_031_d2[7] };
  assign mask_d2_int8_w[32] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20643" *) { vec_data_032_d2[0], vec_data_032_d2[1], vec_data_032_d2[2], vec_data_032_d2[3], vec_data_032_d2[4], vec_data_032_d2[5], vec_data_032_d2[6], vec_data_032_d2[7] };
  assign mask_d2_int8_w[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20644" *) { vec_data_033_d2[0], vec_data_033_d2[1], vec_data_033_d2[2], vec_data_033_d2[3], vec_data_033_d2[4], vec_data_033_d2[5], vec_data_033_d2[6], vec_data_033_d2[7] };
  assign mask_d2_int8_w[34] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20645" *) { vec_data_034_d2[0], vec_data_034_d2[1], vec_data_034_d2[2], vec_data_034_d2[3], vec_data_034_d2[4], vec_data_034_d2[5], vec_data_034_d2[6], vec_data_034_d2[7] };
  assign mask_d2_int8_w[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20646" *) { vec_data_035_d2[0], vec_data_035_d2[1], vec_data_035_d2[2], vec_data_035_d2[3], vec_data_035_d2[4], vec_data_035_d2[5], vec_data_035_d2[6], vec_data_035_d2[7] };
  assign mask_d2_int8_w[36] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20647" *) { vec_data_036_d2[0], vec_data_036_d2[1], vec_data_036_d2[2], vec_data_036_d2[3], vec_data_036_d2[4], vec_data_036_d2[5], vec_data_036_d2[6], vec_data_036_d2[7] };
  assign mask_d2_int8_w[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20648" *) { vec_data_037_d2[0], vec_data_037_d2[1], vec_data_037_d2[2], vec_data_037_d2[3], vec_data_037_d2[4], vec_data_037_d2[5], vec_data_037_d2[6], vec_data_037_d2[7] };
  assign mask_d2_int8_w[38] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20649" *) { vec_data_038_d2[0], vec_data_038_d2[1], vec_data_038_d2[2], vec_data_038_d2[3], vec_data_038_d2[4], vec_data_038_d2[5], vec_data_038_d2[6], vec_data_038_d2[7] };
  assign mask_d2_int8_w[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20650" *) { vec_data_039_d2[0], vec_data_039_d2[1], vec_data_039_d2[2], vec_data_039_d2[3], vec_data_039_d2[4], vec_data_039_d2[5], vec_data_039_d2[6], vec_data_039_d2[7] };
  assign mask_d2_int8_w[40] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20651" *) { vec_data_040_d2[0], vec_data_040_d2[1], vec_data_040_d2[2], vec_data_040_d2[3], vec_data_040_d2[4], vec_data_040_d2[5], vec_data_040_d2[6], vec_data_040_d2[7] };
  assign mask_d2_int8_w[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20652" *) { vec_data_041_d2[0], vec_data_041_d2[1], vec_data_041_d2[2], vec_data_041_d2[3], vec_data_041_d2[4], vec_data_041_d2[5], vec_data_041_d2[6], vec_data_041_d2[7] };
  assign mask_d2_int8_w[42] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20653" *) { vec_data_042_d2[0], vec_data_042_d2[1], vec_data_042_d2[2], vec_data_042_d2[3], vec_data_042_d2[4], vec_data_042_d2[5], vec_data_042_d2[6], vec_data_042_d2[7] };
  assign mask_d2_int8_w[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20654" *) { vec_data_043_d2[0], vec_data_043_d2[1], vec_data_043_d2[2], vec_data_043_d2[3], vec_data_043_d2[4], vec_data_043_d2[5], vec_data_043_d2[6], vec_data_043_d2[7] };
  assign mask_d2_int8_w[44] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20655" *) { vec_data_044_d2[0], vec_data_044_d2[1], vec_data_044_d2[2], vec_data_044_d2[3], vec_data_044_d2[4], vec_data_044_d2[5], vec_data_044_d2[6], vec_data_044_d2[7] };
  assign mask_d2_int8_w[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20656" *) { vec_data_045_d2[0], vec_data_045_d2[1], vec_data_045_d2[2], vec_data_045_d2[3], vec_data_045_d2[4], vec_data_045_d2[5], vec_data_045_d2[6], vec_data_045_d2[7] };
  assign mask_d2_int8_w[46] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20657" *) { vec_data_046_d2[0], vec_data_046_d2[1], vec_data_046_d2[2], vec_data_046_d2[3], vec_data_046_d2[4], vec_data_046_d2[5], vec_data_046_d2[6], vec_data_046_d2[7] };
  assign mask_d2_int8_w[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20658" *) { vec_data_047_d2[0], vec_data_047_d2[1], vec_data_047_d2[2], vec_data_047_d2[3], vec_data_047_d2[4], vec_data_047_d2[5], vec_data_047_d2[6], vec_data_047_d2[7] };
  assign mask_d2_int8_w[48] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20659" *) { vec_data_048_d2[0], vec_data_048_d2[1], vec_data_048_d2[2], vec_data_048_d2[3], vec_data_048_d2[4], vec_data_048_d2[5], vec_data_048_d2[6], vec_data_048_d2[7] };
  assign mask_d2_int8_w[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20660" *) { vec_data_049_d2[0], vec_data_049_d2[1], vec_data_049_d2[2], vec_data_049_d2[3], vec_data_049_d2[4], vec_data_049_d2[5], vec_data_049_d2[6], vec_data_049_d2[7] };
  assign mask_d2_int8_w[50] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20661" *) { vec_data_050_d2[0], vec_data_050_d2[1], vec_data_050_d2[2], vec_data_050_d2[3], vec_data_050_d2[4], vec_data_050_d2[5], vec_data_050_d2[6], vec_data_050_d2[7] };
  assign mask_d2_int8_w[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20662" *) { vec_data_051_d2[0], vec_data_051_d2[1], vec_data_051_d2[2], vec_data_051_d2[3], vec_data_051_d2[4], vec_data_051_d2[5], vec_data_051_d2[6], vec_data_051_d2[7] };
  assign mask_d2_int8_w[52] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20663" *) { vec_data_052_d2[0], vec_data_052_d2[1], vec_data_052_d2[2], vec_data_052_d2[3], vec_data_052_d2[4], vec_data_052_d2[5], vec_data_052_d2[6], vec_data_052_d2[7] };
  assign mask_d2_int8_w[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20664" *) { vec_data_053_d2[0], vec_data_053_d2[1], vec_data_053_d2[2], vec_data_053_d2[3], vec_data_053_d2[4], vec_data_053_d2[5], vec_data_053_d2[6], vec_data_053_d2[7] };
  assign mask_d2_int8_w[54] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20665" *) { vec_data_054_d2[0], vec_data_054_d2[1], vec_data_054_d2[2], vec_data_054_d2[3], vec_data_054_d2[4], vec_data_054_d2[5], vec_data_054_d2[6], vec_data_054_d2[7] };
  assign mask_d2_int8_w[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20666" *) { vec_data_055_d2[0], vec_data_055_d2[1], vec_data_055_d2[2], vec_data_055_d2[3], vec_data_055_d2[4], vec_data_055_d2[5], vec_data_055_d2[6], vec_data_055_d2[7] };
  assign mask_d2_int8_w[56] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20667" *) { vec_data_056_d2[0], vec_data_056_d2[1], vec_data_056_d2[2], vec_data_056_d2[3], vec_data_056_d2[4], vec_data_056_d2[5], vec_data_056_d2[6], vec_data_056_d2[7] };
  assign mask_d2_int8_w[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20668" *) { vec_data_057_d2[0], vec_data_057_d2[1], vec_data_057_d2[2], vec_data_057_d2[3], vec_data_057_d2[4], vec_data_057_d2[5], vec_data_057_d2[6], vec_data_057_d2[7] };
  assign mask_d2_int8_w[58] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20669" *) { vec_data_058_d2[0], vec_data_058_d2[1], vec_data_058_d2[2], vec_data_058_d2[3], vec_data_058_d2[4], vec_data_058_d2[5], vec_data_058_d2[6], vec_data_058_d2[7] };
  assign mask_d2_int8_w[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20670" *) { vec_data_059_d2[0], vec_data_059_d2[1], vec_data_059_d2[2], vec_data_059_d2[3], vec_data_059_d2[4], vec_data_059_d2[5], vec_data_059_d2[6], vec_data_059_d2[7] };
  assign mask_d2_int8_w[60] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20671" *) { vec_data_060_d2[0], vec_data_060_d2[1], vec_data_060_d2[2], vec_data_060_d2[3], vec_data_060_d2[4], vec_data_060_d2[5], vec_data_060_d2[6], vec_data_060_d2[7] };
  assign mask_d2_int8_w[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20672" *) { vec_data_061_d2[0], vec_data_061_d2[1], vec_data_061_d2[2], vec_data_061_d2[3], vec_data_061_d2[4], vec_data_061_d2[5], vec_data_061_d2[6], vec_data_061_d2[7] };
  assign mask_d2_int8_w[62] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20673" *) { vec_data_062_d2[0], vec_data_062_d2[1], vec_data_062_d2[2], vec_data_062_d2[3], vec_data_062_d2[4], vec_data_062_d2[5], vec_data_062_d2[6], vec_data_062_d2[7] };
  assign mask_d2_int8_w[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20674" *) { vec_data_063_d2[0], vec_data_063_d2[1], vec_data_063_d2[2], vec_data_063_d2[3], vec_data_063_d2[4], vec_data_063_d2[5], vec_data_063_d2[6], vec_data_063_d2[7] };
  assign mask_d2_int8_w[64] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20675" *) { vec_data_064_d2[0], vec_data_064_d2[1], vec_data_064_d2[2], vec_data_064_d2[3], vec_data_064_d2[4], vec_data_064_d2[5], vec_data_064_d2[6], vec_data_064_d2[7] };
  assign mask_d2_int8_w[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20676" *) { vec_data_065_d2[0], vec_data_065_d2[1], vec_data_065_d2[2], vec_data_065_d2[3], vec_data_065_d2[4], vec_data_065_d2[5], vec_data_065_d2[6], vec_data_065_d2[7] };
  assign mask_d2_int8_w[66] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20677" *) { vec_data_066_d2[0], vec_data_066_d2[1], vec_data_066_d2[2], vec_data_066_d2[3], vec_data_066_d2[4], vec_data_066_d2[5], vec_data_066_d2[6], vec_data_066_d2[7] };
  assign mask_d2_int8_w[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20678" *) { vec_data_067_d2[0], vec_data_067_d2[1], vec_data_067_d2[2], vec_data_067_d2[3], vec_data_067_d2[4], vec_data_067_d2[5], vec_data_067_d2[6], vec_data_067_d2[7] };
  assign mask_d2_int8_w[68] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20679" *) { vec_data_068_d2[0], vec_data_068_d2[1], vec_data_068_d2[2], vec_data_068_d2[3], vec_data_068_d2[4], vec_data_068_d2[5], vec_data_068_d2[6], vec_data_068_d2[7] };
  assign mask_d2_int8_w[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20680" *) { vec_data_069_d2[0], vec_data_069_d2[1], vec_data_069_d2[2], vec_data_069_d2[3], vec_data_069_d2[4], vec_data_069_d2[5], vec_data_069_d2[6], vec_data_069_d2[7] };
  assign mask_d2_int8_w[70] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20681" *) { vec_data_070_d2[0], vec_data_070_d2[1], vec_data_070_d2[2], vec_data_070_d2[3], vec_data_070_d2[4], vec_data_070_d2[5], vec_data_070_d2[6], vec_data_070_d2[7] };
  assign mask_d2_int8_w[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20682" *) { vec_data_071_d2[0], vec_data_071_d2[1], vec_data_071_d2[2], vec_data_071_d2[3], vec_data_071_d2[4], vec_data_071_d2[5], vec_data_071_d2[6], vec_data_071_d2[7] };
  assign mask_d2_int8_w[72] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20683" *) { vec_data_072_d2[0], vec_data_072_d2[1], vec_data_072_d2[2], vec_data_072_d2[3], vec_data_072_d2[4], vec_data_072_d2[5], vec_data_072_d2[6], vec_data_072_d2[7] };
  assign mask_d2_int8_w[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20684" *) { vec_data_073_d2[0], vec_data_073_d2[1], vec_data_073_d2[2], vec_data_073_d2[3], vec_data_073_d2[4], vec_data_073_d2[5], vec_data_073_d2[6], vec_data_073_d2[7] };
  assign mask_d2_int8_w[74] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20685" *) { vec_data_074_d2[0], vec_data_074_d2[1], vec_data_074_d2[2], vec_data_074_d2[3], vec_data_074_d2[4], vec_data_074_d2[5], vec_data_074_d2[6], vec_data_074_d2[7] };
  assign mask_d2_int8_w[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20686" *) { vec_data_075_d2[0], vec_data_075_d2[1], vec_data_075_d2[2], vec_data_075_d2[3], vec_data_075_d2[4], vec_data_075_d2[5], vec_data_075_d2[6], vec_data_075_d2[7] };
  assign mask_d2_int8_w[76] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20687" *) { vec_data_076_d2[0], vec_data_076_d2[1], vec_data_076_d2[2], vec_data_076_d2[3], vec_data_076_d2[4], vec_data_076_d2[5], vec_data_076_d2[6], vec_data_076_d2[7] };
  assign mask_d2_int8_w[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20688" *) { vec_data_077_d2[0], vec_data_077_d2[1], vec_data_077_d2[2], vec_data_077_d2[3], vec_data_077_d2[4], vec_data_077_d2[5], vec_data_077_d2[6], vec_data_077_d2[7] };
  assign mask_d2_int8_w[78] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20689" *) { vec_data_078_d2[0], vec_data_078_d2[1], vec_data_078_d2[2], vec_data_078_d2[3], vec_data_078_d2[4], vec_data_078_d2[5], vec_data_078_d2[6], vec_data_078_d2[7] };
  assign mask_d2_int8_w[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20690" *) { vec_data_079_d2[0], vec_data_079_d2[1], vec_data_079_d2[2], vec_data_079_d2[3], vec_data_079_d2[4], vec_data_079_d2[5], vec_data_079_d2[6], vec_data_079_d2[7] };
  assign mask_d2_int8_w[80] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20691" *) { vec_data_080_d2[0], vec_data_080_d2[1], vec_data_080_d2[2], vec_data_080_d2[3], vec_data_080_d2[4], vec_data_080_d2[5], vec_data_080_d2[6], vec_data_080_d2[7] };
  assign mask_d2_int8_w[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20692" *) { vec_data_081_d2[0], vec_data_081_d2[1], vec_data_081_d2[2], vec_data_081_d2[3], vec_data_081_d2[4], vec_data_081_d2[5], vec_data_081_d2[6], vec_data_081_d2[7] };
  assign mask_d2_int8_w[82] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20693" *) { vec_data_082_d2[0], vec_data_082_d2[1], vec_data_082_d2[2], vec_data_082_d2[3], vec_data_082_d2[4], vec_data_082_d2[5], vec_data_082_d2[6], vec_data_082_d2[7] };
  assign mask_d2_int8_w[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20694" *) { vec_data_083_d2[0], vec_data_083_d2[1], vec_data_083_d2[2], vec_data_083_d2[3], vec_data_083_d2[4], vec_data_083_d2[5], vec_data_083_d2[6], vec_data_083_d2[7] };
  assign mask_d2_int8_w[84] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20695" *) { vec_data_084_d2[0], vec_data_084_d2[1], vec_data_084_d2[2], vec_data_084_d2[3], vec_data_084_d2[4], vec_data_084_d2[5], vec_data_084_d2[6], vec_data_084_d2[7] };
  assign mask_d2_int8_w[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20696" *) { vec_data_085_d2[0], vec_data_085_d2[1], vec_data_085_d2[2], vec_data_085_d2[3], vec_data_085_d2[4], vec_data_085_d2[5], vec_data_085_d2[6], vec_data_085_d2[7] };
  assign mask_d2_int8_w[86] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20697" *) { vec_data_086_d2[0], vec_data_086_d2[1], vec_data_086_d2[2], vec_data_086_d2[3], vec_data_086_d2[4], vec_data_086_d2[5], vec_data_086_d2[6], vec_data_086_d2[7] };
  assign mask_d2_int8_w[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20698" *) { vec_data_087_d2[0], vec_data_087_d2[1], vec_data_087_d2[2], vec_data_087_d2[3], vec_data_087_d2[4], vec_data_087_d2[5], vec_data_087_d2[6], vec_data_087_d2[7] };
  assign mask_d2_int8_w[88] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20699" *) { vec_data_088_d2[0], vec_data_088_d2[1], vec_data_088_d2[2], vec_data_088_d2[3], vec_data_088_d2[4], vec_data_088_d2[5], vec_data_088_d2[6], vec_data_088_d2[7] };
  assign mask_d2_int8_w[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20700" *) { vec_data_089_d2[0], vec_data_089_d2[1], vec_data_089_d2[2], vec_data_089_d2[3], vec_data_089_d2[4], vec_data_089_d2[5], vec_data_089_d2[6], vec_data_089_d2[7] };
  assign mask_d2_int8_w[90] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20701" *) { vec_data_090_d2[0], vec_data_090_d2[1], vec_data_090_d2[2], vec_data_090_d2[3], vec_data_090_d2[4], vec_data_090_d2[5], vec_data_090_d2[6], vec_data_090_d2[7] };
  assign mask_d2_int8_w[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20702" *) { vec_data_091_d2[0], vec_data_091_d2[1], vec_data_091_d2[2], vec_data_091_d2[3], vec_data_091_d2[4], vec_data_091_d2[5], vec_data_091_d2[6], vec_data_091_d2[7] };
  assign mask_d2_int8_w[92] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20703" *) { vec_data_092_d2[0], vec_data_092_d2[1], vec_data_092_d2[2], vec_data_092_d2[3], vec_data_092_d2[4], vec_data_092_d2[5], vec_data_092_d2[6], vec_data_092_d2[7] };
  assign mask_d2_int8_w[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20704" *) { vec_data_093_d2[0], vec_data_093_d2[1], vec_data_093_d2[2], vec_data_093_d2[3], vec_data_093_d2[4], vec_data_093_d2[5], vec_data_093_d2[6], vec_data_093_d2[7] };
  assign mask_d2_int8_w[94] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20705" *) { vec_data_094_d2[0], vec_data_094_d2[1], vec_data_094_d2[2], vec_data_094_d2[3], vec_data_094_d2[4], vec_data_094_d2[5], vec_data_094_d2[6], vec_data_094_d2[7] };
  assign mask_d2_int8_w[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20706" *) { vec_data_095_d2[0], vec_data_095_d2[1], vec_data_095_d2[2], vec_data_095_d2[3], vec_data_095_d2[4], vec_data_095_d2[5], vec_data_095_d2[6], vec_data_095_d2[7] };
  assign mask_d2_int8_w[96] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20707" *) { vec_data_096_d2[0], vec_data_096_d2[1], vec_data_096_d2[2], vec_data_096_d2[3], vec_data_096_d2[4], vec_data_096_d2[5], vec_data_096_d2[6], vec_data_096_d2[7] };
  assign mask_d2_int8_w[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20708" *) { vec_data_097_d2[0], vec_data_097_d2[1], vec_data_097_d2[2], vec_data_097_d2[3], vec_data_097_d2[4], vec_data_097_d2[5], vec_data_097_d2[6], vec_data_097_d2[7] };
  assign mask_d2_int8_w[98] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20709" *) { vec_data_098_d2[0], vec_data_098_d2[1], vec_data_098_d2[2], vec_data_098_d2[3], vec_data_098_d2[4], vec_data_098_d2[5], vec_data_098_d2[6], vec_data_098_d2[7] };
  assign mask_d2_int8_w[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20710" *) { vec_data_099_d2[0], vec_data_099_d2[1], vec_data_099_d2[2], vec_data_099_d2[3], vec_data_099_d2[4], vec_data_099_d2[5], vec_data_099_d2[6], vec_data_099_d2[7] };
  assign mask_d2_int8_w[100] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20711" *) { vec_data_100_d2[0], vec_data_100_d2[1], vec_data_100_d2[2], vec_data_100_d2[3], vec_data_100_d2[4], vec_data_100_d2[5], vec_data_100_d2[6], vec_data_100_d2[7] };
  assign mask_d2_int8_w[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20712" *) { vec_data_101_d2[0], vec_data_101_d2[1], vec_data_101_d2[2], vec_data_101_d2[3], vec_data_101_d2[4], vec_data_101_d2[5], vec_data_101_d2[6], vec_data_101_d2[7] };
  assign mask_d2_int8_w[102] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20713" *) { vec_data_102_d2[0], vec_data_102_d2[1], vec_data_102_d2[2], vec_data_102_d2[3], vec_data_102_d2[4], vec_data_102_d2[5], vec_data_102_d2[6], vec_data_102_d2[7] };
  assign mask_d2_int8_w[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20714" *) { vec_data_103_d2[0], vec_data_103_d2[1], vec_data_103_d2[2], vec_data_103_d2[3], vec_data_103_d2[4], vec_data_103_d2[5], vec_data_103_d2[6], vec_data_103_d2[7] };
  assign mask_d2_int8_w[104] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20715" *) { vec_data_104_d2[0], vec_data_104_d2[1], vec_data_104_d2[2], vec_data_104_d2[3], vec_data_104_d2[4], vec_data_104_d2[5], vec_data_104_d2[6], vec_data_104_d2[7] };
  assign mask_d2_int8_w[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20716" *) { vec_data_105_d2[0], vec_data_105_d2[1], vec_data_105_d2[2], vec_data_105_d2[3], vec_data_105_d2[4], vec_data_105_d2[5], vec_data_105_d2[6], vec_data_105_d2[7] };
  assign mask_d2_int8_w[106] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20717" *) { vec_data_106_d2[0], vec_data_106_d2[1], vec_data_106_d2[2], vec_data_106_d2[3], vec_data_106_d2[4], vec_data_106_d2[5], vec_data_106_d2[6], vec_data_106_d2[7] };
  assign mask_d2_int8_w[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20718" *) { vec_data_107_d2[0], vec_data_107_d2[1], vec_data_107_d2[2], vec_data_107_d2[3], vec_data_107_d2[4], vec_data_107_d2[5], vec_data_107_d2[6], vec_data_107_d2[7] };
  assign mask_d2_int8_w[108] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20719" *) { vec_data_108_d2[0], vec_data_108_d2[1], vec_data_108_d2[2], vec_data_108_d2[3], vec_data_108_d2[4], vec_data_108_d2[5], vec_data_108_d2[6], vec_data_108_d2[7] };
  assign mask_d2_int8_w[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20720" *) { vec_data_109_d2[0], vec_data_109_d2[1], vec_data_109_d2[2], vec_data_109_d2[3], vec_data_109_d2[4], vec_data_109_d2[5], vec_data_109_d2[6], vec_data_109_d2[7] };
  assign mask_d2_int8_w[110] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20721" *) { vec_data_110_d2[0], vec_data_110_d2[1], vec_data_110_d2[2], vec_data_110_d2[3], vec_data_110_d2[4], vec_data_110_d2[5], vec_data_110_d2[6], vec_data_110_d2[7] };
  assign mask_d2_int8_w[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20722" *) { vec_data_111_d2[0], vec_data_111_d2[1], vec_data_111_d2[2], vec_data_111_d2[3], vec_data_111_d2[4], vec_data_111_d2[5], vec_data_111_d2[6], vec_data_111_d2[7] };
  assign mask_d2_int8_w[112] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20723" *) { vec_data_112_d2[0], vec_data_112_d2[1], vec_data_112_d2[2], vec_data_112_d2[3], vec_data_112_d2[4], vec_data_112_d2[5], vec_data_112_d2[6], vec_data_112_d2[7] };
  assign mask_d2_int8_w[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20724" *) { vec_data_113_d2[0], vec_data_113_d2[1], vec_data_113_d2[2], vec_data_113_d2[3], vec_data_113_d2[4], vec_data_113_d2[5], vec_data_113_d2[6], vec_data_113_d2[7] };
  assign mask_d2_int8_w[114] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20725" *) { vec_data_114_d2[0], vec_data_114_d2[1], vec_data_114_d2[2], vec_data_114_d2[3], vec_data_114_d2[4], vec_data_114_d2[5], vec_data_114_d2[6], vec_data_114_d2[7] };
  assign mask_d2_int8_w[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20726" *) { vec_data_115_d2[0], vec_data_115_d2[1], vec_data_115_d2[2], vec_data_115_d2[3], vec_data_115_d2[4], vec_data_115_d2[5], vec_data_115_d2[6], vec_data_115_d2[7] };
  assign mask_d2_int8_w[116] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20727" *) { vec_data_116_d2[0], vec_data_116_d2[1], vec_data_116_d2[2], vec_data_116_d2[3], vec_data_116_d2[4], vec_data_116_d2[5], vec_data_116_d2[6], vec_data_116_d2[7] };
  assign mask_d2_int8_w[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20728" *) { vec_data_117_d2[0], vec_data_117_d2[1], vec_data_117_d2[2], vec_data_117_d2[3], vec_data_117_d2[4], vec_data_117_d2[5], vec_data_117_d2[6], vec_data_117_d2[7] };
  assign mask_d2_int8_w[118] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20729" *) { vec_data_118_d2[0], vec_data_118_d2[1], vec_data_118_d2[2], vec_data_118_d2[3], vec_data_118_d2[4], vec_data_118_d2[5], vec_data_118_d2[6], vec_data_118_d2[7] };
  assign mask_d2_int8_w[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20730" *) { vec_data_119_d2[0], vec_data_119_d2[1], vec_data_119_d2[2], vec_data_119_d2[3], vec_data_119_d2[4], vec_data_119_d2[5], vec_data_119_d2[6], vec_data_119_d2[7] };
  assign mask_d2_int8_w[120] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20731" *) { vec_data_120_d2[0], vec_data_120_d2[1], vec_data_120_d2[2], vec_data_120_d2[3], vec_data_120_d2[4], vec_data_120_d2[5], vec_data_120_d2[6], vec_data_120_d2[7] };
  assign mask_d2_int8_w[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20732" *) { vec_data_121_d2[0], vec_data_121_d2[1], vec_data_121_d2[2], vec_data_121_d2[3], vec_data_121_d2[4], vec_data_121_d2[5], vec_data_121_d2[6], vec_data_121_d2[7] };
  assign mask_d2_int8_w[122] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20733" *) { vec_data_122_d2[0], vec_data_122_d2[1], vec_data_122_d2[2], vec_data_122_d2[3], vec_data_122_d2[4], vec_data_122_d2[5], vec_data_122_d2[6], vec_data_122_d2[7] };
  assign mask_d2_int8_w[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20734" *) { vec_data_123_d2[0], vec_data_123_d2[1], vec_data_123_d2[2], vec_data_123_d2[3], vec_data_123_d2[4], vec_data_123_d2[5], vec_data_123_d2[6], vec_data_123_d2[7] };
  assign mask_d2_int8_w[124] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20735" *) { vec_data_124_d2[0], vec_data_124_d2[1], vec_data_124_d2[2], vec_data_124_d2[3], vec_data_124_d2[4], vec_data_124_d2[5], vec_data_124_d2[6], vec_data_124_d2[7] };
  assign mask_d2_int8_w[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20736" *) { vec_data_125_d2[0], vec_data_125_d2[1], vec_data_125_d2[2], vec_data_125_d2[3], vec_data_125_d2[4], vec_data_125_d2[5], vec_data_125_d2[6], vec_data_125_d2[7] };
  assign mask_d2_int8_w[126] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20737" *) { vec_data_126_d2[0], vec_data_126_d2[1], vec_data_126_d2[2], vec_data_126_d2[3], vec_data_126_d2[4], vec_data_126_d2[5], vec_data_126_d2[6], vec_data_126_d2[7] };
  assign mask_d2_int8_w[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20738" *) { vec_data_127_d2[0], vec_data_127_d2[1], vec_data_127_d2[2], vec_data_127_d2[3], vec_data_127_d2[4], vec_data_127_d2[5], vec_data_127_d2[6], vec_data_127_d2[7] };
  assign mask_d2_int16_w[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20870" *) { vec_data_000_d2[0], vec_data_000_d2[1], vec_data_000_d2[2], vec_data_000_d2[3], vec_data_000_d2[4], vec_data_000_d2[5], vec_data_000_d2[6], vec_data_000_d2[7], vec_data_001_d2[0], vec_data_001_d2[1], vec_data_001_d2[2], vec_data_001_d2[3], vec_data_001_d2[4], vec_data_001_d2[5], vec_data_001_d2[6], vec_data_001_d2[7] };
  assign mask_d2_int16_w[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20871" *) { vec_data_002_d2[0], vec_data_002_d2[1], vec_data_002_d2[2], vec_data_002_d2[3], vec_data_002_d2[4], vec_data_002_d2[5], vec_data_002_d2[6], vec_data_002_d2[7], vec_data_003_d2[0], vec_data_003_d2[1], vec_data_003_d2[2], vec_data_003_d2[3], vec_data_003_d2[4], vec_data_003_d2[5], vec_data_003_d2[6], vec_data_003_d2[7] };
  assign mask_d2_int16_w[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20872" *) { vec_data_004_d2[0], vec_data_004_d2[1], vec_data_004_d2[2], vec_data_004_d2[3], vec_data_004_d2[4], vec_data_004_d2[5], vec_data_004_d2[6], vec_data_004_d2[7], vec_data_005_d2[0], vec_data_005_d2[1], vec_data_005_d2[2], vec_data_005_d2[3], vec_data_005_d2[4], vec_data_005_d2[5], vec_data_005_d2[6], vec_data_005_d2[7] };
  assign mask_d2_int16_w[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20873" *) { vec_data_006_d2[0], vec_data_006_d2[1], vec_data_006_d2[2], vec_data_006_d2[3], vec_data_006_d2[4], vec_data_006_d2[5], vec_data_006_d2[6], vec_data_006_d2[7], vec_data_007_d2[0], vec_data_007_d2[1], vec_data_007_d2[2], vec_data_007_d2[3], vec_data_007_d2[4], vec_data_007_d2[5], vec_data_007_d2[6], vec_data_007_d2[7] };
  assign mask_d2_int16_w[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20874" *) { vec_data_008_d2[0], vec_data_008_d2[1], vec_data_008_d2[2], vec_data_008_d2[3], vec_data_008_d2[4], vec_data_008_d2[5], vec_data_008_d2[6], vec_data_008_d2[7], vec_data_009_d2[0], vec_data_009_d2[1], vec_data_009_d2[2], vec_data_009_d2[3], vec_data_009_d2[4], vec_data_009_d2[5], vec_data_009_d2[6], vec_data_009_d2[7] };
  assign mask_d2_int16_w[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20875" *) { vec_data_010_d2[0], vec_data_010_d2[1], vec_data_010_d2[2], vec_data_010_d2[3], vec_data_010_d2[4], vec_data_010_d2[5], vec_data_010_d2[6], vec_data_010_d2[7], vec_data_011_d2[0], vec_data_011_d2[1], vec_data_011_d2[2], vec_data_011_d2[3], vec_data_011_d2[4], vec_data_011_d2[5], vec_data_011_d2[6], vec_data_011_d2[7] };
  assign mask_d2_int16_w[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20876" *) { vec_data_012_d2[0], vec_data_012_d2[1], vec_data_012_d2[2], vec_data_012_d2[3], vec_data_012_d2[4], vec_data_012_d2[5], vec_data_012_d2[6], vec_data_012_d2[7], vec_data_013_d2[0], vec_data_013_d2[1], vec_data_013_d2[2], vec_data_013_d2[3], vec_data_013_d2[4], vec_data_013_d2[5], vec_data_013_d2[6], vec_data_013_d2[7] };
  assign mask_d2_int16_w[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20877" *) { vec_data_014_d2[0], vec_data_014_d2[1], vec_data_014_d2[2], vec_data_014_d2[3], vec_data_014_d2[4], vec_data_014_d2[5], vec_data_014_d2[6], vec_data_014_d2[7], vec_data_015_d2[0], vec_data_015_d2[1], vec_data_015_d2[2], vec_data_015_d2[3], vec_data_015_d2[4], vec_data_015_d2[5], vec_data_015_d2[6], vec_data_015_d2[7] };
  assign mask_d2_int16_w[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20878" *) { vec_data_016_d2[0], vec_data_016_d2[1], vec_data_016_d2[2], vec_data_016_d2[3], vec_data_016_d2[4], vec_data_016_d2[5], vec_data_016_d2[6], vec_data_016_d2[7], vec_data_017_d2[0], vec_data_017_d2[1], vec_data_017_d2[2], vec_data_017_d2[3], vec_data_017_d2[4], vec_data_017_d2[5], vec_data_017_d2[6], vec_data_017_d2[7] };
  assign mask_d2_int16_w[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20879" *) { vec_data_018_d2[0], vec_data_018_d2[1], vec_data_018_d2[2], vec_data_018_d2[3], vec_data_018_d2[4], vec_data_018_d2[5], vec_data_018_d2[6], vec_data_018_d2[7], vec_data_019_d2[0], vec_data_019_d2[1], vec_data_019_d2[2], vec_data_019_d2[3], vec_data_019_d2[4], vec_data_019_d2[5], vec_data_019_d2[6], vec_data_019_d2[7] };
  assign mask_d2_int16_w[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20880" *) { vec_data_020_d2[0], vec_data_020_d2[1], vec_data_020_d2[2], vec_data_020_d2[3], vec_data_020_d2[4], vec_data_020_d2[5], vec_data_020_d2[6], vec_data_020_d2[7], vec_data_021_d2[0], vec_data_021_d2[1], vec_data_021_d2[2], vec_data_021_d2[3], vec_data_021_d2[4], vec_data_021_d2[5], vec_data_021_d2[6], vec_data_021_d2[7] };
  assign mask_d2_int16_w[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20881" *) { vec_data_022_d2[0], vec_data_022_d2[1], vec_data_022_d2[2], vec_data_022_d2[3], vec_data_022_d2[4], vec_data_022_d2[5], vec_data_022_d2[6], vec_data_022_d2[7], vec_data_023_d2[0], vec_data_023_d2[1], vec_data_023_d2[2], vec_data_023_d2[3], vec_data_023_d2[4], vec_data_023_d2[5], vec_data_023_d2[6], vec_data_023_d2[7] };
  assign mask_d2_int16_w[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20882" *) { vec_data_024_d2[0], vec_data_024_d2[1], vec_data_024_d2[2], vec_data_024_d2[3], vec_data_024_d2[4], vec_data_024_d2[5], vec_data_024_d2[6], vec_data_024_d2[7], vec_data_025_d2[0], vec_data_025_d2[1], vec_data_025_d2[2], vec_data_025_d2[3], vec_data_025_d2[4], vec_data_025_d2[5], vec_data_025_d2[6], vec_data_025_d2[7] };
  assign mask_d2_int16_w[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20883" *) { vec_data_026_d2[0], vec_data_026_d2[1], vec_data_026_d2[2], vec_data_026_d2[3], vec_data_026_d2[4], vec_data_026_d2[5], vec_data_026_d2[6], vec_data_026_d2[7], vec_data_027_d2[0], vec_data_027_d2[1], vec_data_027_d2[2], vec_data_027_d2[3], vec_data_027_d2[4], vec_data_027_d2[5], vec_data_027_d2[6], vec_data_027_d2[7] };
  assign mask_d2_int16_w[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20884" *) { vec_data_028_d2[0], vec_data_028_d2[1], vec_data_028_d2[2], vec_data_028_d2[3], vec_data_028_d2[4], vec_data_028_d2[5], vec_data_028_d2[6], vec_data_028_d2[7], vec_data_029_d2[0], vec_data_029_d2[1], vec_data_029_d2[2], vec_data_029_d2[3], vec_data_029_d2[4], vec_data_029_d2[5], vec_data_029_d2[6], vec_data_029_d2[7] };
  assign mask_d2_int16_w[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20885" *) { vec_data_030_d2[0], vec_data_030_d2[1], vec_data_030_d2[2], vec_data_030_d2[3], vec_data_030_d2[4], vec_data_030_d2[5], vec_data_030_d2[6], vec_data_030_d2[7], vec_data_031_d2[0], vec_data_031_d2[1], vec_data_031_d2[2], vec_data_031_d2[3], vec_data_031_d2[4], vec_data_031_d2[5], vec_data_031_d2[6], vec_data_031_d2[7] };
  assign mask_d2_int16_w[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20886" *) { vec_data_032_d2[0], vec_data_032_d2[1], vec_data_032_d2[2], vec_data_032_d2[3], vec_data_032_d2[4], vec_data_032_d2[5], vec_data_032_d2[6], vec_data_032_d2[7], vec_data_033_d2[0], vec_data_033_d2[1], vec_data_033_d2[2], vec_data_033_d2[3], vec_data_033_d2[4], vec_data_033_d2[5], vec_data_033_d2[6], vec_data_033_d2[7] };
  assign mask_d2_int16_w[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20887" *) { vec_data_034_d2[0], vec_data_034_d2[1], vec_data_034_d2[2], vec_data_034_d2[3], vec_data_034_d2[4], vec_data_034_d2[5], vec_data_034_d2[6], vec_data_034_d2[7], vec_data_035_d2[0], vec_data_035_d2[1], vec_data_035_d2[2], vec_data_035_d2[3], vec_data_035_d2[4], vec_data_035_d2[5], vec_data_035_d2[6], vec_data_035_d2[7] };
  assign mask_d2_int16_w[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20888" *) { vec_data_036_d2[0], vec_data_036_d2[1], vec_data_036_d2[2], vec_data_036_d2[3], vec_data_036_d2[4], vec_data_036_d2[5], vec_data_036_d2[6], vec_data_036_d2[7], vec_data_037_d2[0], vec_data_037_d2[1], vec_data_037_d2[2], vec_data_037_d2[3], vec_data_037_d2[4], vec_data_037_d2[5], vec_data_037_d2[6], vec_data_037_d2[7] };
  assign mask_d2_int16_w[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20889" *) { vec_data_038_d2[0], vec_data_038_d2[1], vec_data_038_d2[2], vec_data_038_d2[3], vec_data_038_d2[4], vec_data_038_d2[5], vec_data_038_d2[6], vec_data_038_d2[7], vec_data_039_d2[0], vec_data_039_d2[1], vec_data_039_d2[2], vec_data_039_d2[3], vec_data_039_d2[4], vec_data_039_d2[5], vec_data_039_d2[6], vec_data_039_d2[7] };
  assign mask_d2_int16_w[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20890" *) { vec_data_040_d2[0], vec_data_040_d2[1], vec_data_040_d2[2], vec_data_040_d2[3], vec_data_040_d2[4], vec_data_040_d2[5], vec_data_040_d2[6], vec_data_040_d2[7], vec_data_041_d2[0], vec_data_041_d2[1], vec_data_041_d2[2], vec_data_041_d2[3], vec_data_041_d2[4], vec_data_041_d2[5], vec_data_041_d2[6], vec_data_041_d2[7] };
  assign mask_d2_int16_w[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20891" *) { vec_data_042_d2[0], vec_data_042_d2[1], vec_data_042_d2[2], vec_data_042_d2[3], vec_data_042_d2[4], vec_data_042_d2[5], vec_data_042_d2[6], vec_data_042_d2[7], vec_data_043_d2[0], vec_data_043_d2[1], vec_data_043_d2[2], vec_data_043_d2[3], vec_data_043_d2[4], vec_data_043_d2[5], vec_data_043_d2[6], vec_data_043_d2[7] };
  assign mask_d2_int16_w[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20892" *) { vec_data_044_d2[0], vec_data_044_d2[1], vec_data_044_d2[2], vec_data_044_d2[3], vec_data_044_d2[4], vec_data_044_d2[5], vec_data_044_d2[6], vec_data_044_d2[7], vec_data_045_d2[0], vec_data_045_d2[1], vec_data_045_d2[2], vec_data_045_d2[3], vec_data_045_d2[4], vec_data_045_d2[5], vec_data_045_d2[6], vec_data_045_d2[7] };
  assign mask_d2_int16_w[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20893" *) { vec_data_046_d2[0], vec_data_046_d2[1], vec_data_046_d2[2], vec_data_046_d2[3], vec_data_046_d2[4], vec_data_046_d2[5], vec_data_046_d2[6], vec_data_046_d2[7], vec_data_047_d2[0], vec_data_047_d2[1], vec_data_047_d2[2], vec_data_047_d2[3], vec_data_047_d2[4], vec_data_047_d2[5], vec_data_047_d2[6], vec_data_047_d2[7] };
  assign mask_d2_int16_w[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20894" *) { vec_data_048_d2[0], vec_data_048_d2[1], vec_data_048_d2[2], vec_data_048_d2[3], vec_data_048_d2[4], vec_data_048_d2[5], vec_data_048_d2[6], vec_data_048_d2[7], vec_data_049_d2[0], vec_data_049_d2[1], vec_data_049_d2[2], vec_data_049_d2[3], vec_data_049_d2[4], vec_data_049_d2[5], vec_data_049_d2[6], vec_data_049_d2[7] };
  assign mask_d2_int16_w[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20895" *) { vec_data_050_d2[0], vec_data_050_d2[1], vec_data_050_d2[2], vec_data_050_d2[3], vec_data_050_d2[4], vec_data_050_d2[5], vec_data_050_d2[6], vec_data_050_d2[7], vec_data_051_d2[0], vec_data_051_d2[1], vec_data_051_d2[2], vec_data_051_d2[3], vec_data_051_d2[4], vec_data_051_d2[5], vec_data_051_d2[6], vec_data_051_d2[7] };
  assign mask_d2_int16_w[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20896" *) { vec_data_052_d2[0], vec_data_052_d2[1], vec_data_052_d2[2], vec_data_052_d2[3], vec_data_052_d2[4], vec_data_052_d2[5], vec_data_052_d2[6], vec_data_052_d2[7], vec_data_053_d2[0], vec_data_053_d2[1], vec_data_053_d2[2], vec_data_053_d2[3], vec_data_053_d2[4], vec_data_053_d2[5], vec_data_053_d2[6], vec_data_053_d2[7] };
  assign mask_d2_int16_w[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20897" *) { vec_data_054_d2[0], vec_data_054_d2[1], vec_data_054_d2[2], vec_data_054_d2[3], vec_data_054_d2[4], vec_data_054_d2[5], vec_data_054_d2[6], vec_data_054_d2[7], vec_data_055_d2[0], vec_data_055_d2[1], vec_data_055_d2[2], vec_data_055_d2[3], vec_data_055_d2[4], vec_data_055_d2[5], vec_data_055_d2[6], vec_data_055_d2[7] };
  assign mask_d2_int16_w[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20898" *) { vec_data_056_d2[0], vec_data_056_d2[1], vec_data_056_d2[2], vec_data_056_d2[3], vec_data_056_d2[4], vec_data_056_d2[5], vec_data_056_d2[6], vec_data_056_d2[7], vec_data_057_d2[0], vec_data_057_d2[1], vec_data_057_d2[2], vec_data_057_d2[3], vec_data_057_d2[4], vec_data_057_d2[5], vec_data_057_d2[6], vec_data_057_d2[7] };
  assign mask_d2_int16_w[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20899" *) { vec_data_058_d2[0], vec_data_058_d2[1], vec_data_058_d2[2], vec_data_058_d2[3], vec_data_058_d2[4], vec_data_058_d2[5], vec_data_058_d2[6], vec_data_058_d2[7], vec_data_059_d2[0], vec_data_059_d2[1], vec_data_059_d2[2], vec_data_059_d2[3], vec_data_059_d2[4], vec_data_059_d2[5], vec_data_059_d2[6], vec_data_059_d2[7] };
  assign mask_d2_int16_w[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20900" *) { vec_data_060_d2[0], vec_data_060_d2[1], vec_data_060_d2[2], vec_data_060_d2[3], vec_data_060_d2[4], vec_data_060_d2[5], vec_data_060_d2[6], vec_data_060_d2[7], vec_data_061_d2[0], vec_data_061_d2[1], vec_data_061_d2[2], vec_data_061_d2[3], vec_data_061_d2[4], vec_data_061_d2[5], vec_data_061_d2[6], vec_data_061_d2[7] };
  assign mask_d2_int16_w[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20901" *) { vec_data_062_d2[0], vec_data_062_d2[1], vec_data_062_d2[2], vec_data_062_d2[3], vec_data_062_d2[4], vec_data_062_d2[5], vec_data_062_d2[6], vec_data_062_d2[7], vec_data_063_d2[0], vec_data_063_d2[1], vec_data_063_d2[2], vec_data_063_d2[3], vec_data_063_d2[4], vec_data_063_d2[5], vec_data_063_d2[6], vec_data_063_d2[7] };
  assign mask_d2_int16_w[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20902" *) { vec_data_064_d2[0], vec_data_064_d2[1], vec_data_064_d2[2], vec_data_064_d2[3], vec_data_064_d2[4], vec_data_064_d2[5], vec_data_064_d2[6], vec_data_064_d2[7], vec_data_065_d2[0], vec_data_065_d2[1], vec_data_065_d2[2], vec_data_065_d2[3], vec_data_065_d2[4], vec_data_065_d2[5], vec_data_065_d2[6], vec_data_065_d2[7] };
  assign mask_d2_int16_w[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20903" *) { vec_data_066_d2[0], vec_data_066_d2[1], vec_data_066_d2[2], vec_data_066_d2[3], vec_data_066_d2[4], vec_data_066_d2[5], vec_data_066_d2[6], vec_data_066_d2[7], vec_data_067_d2[0], vec_data_067_d2[1], vec_data_067_d2[2], vec_data_067_d2[3], vec_data_067_d2[4], vec_data_067_d2[5], vec_data_067_d2[6], vec_data_067_d2[7] };
  assign mask_d2_int16_w[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20904" *) { vec_data_068_d2[0], vec_data_068_d2[1], vec_data_068_d2[2], vec_data_068_d2[3], vec_data_068_d2[4], vec_data_068_d2[5], vec_data_068_d2[6], vec_data_068_d2[7], vec_data_069_d2[0], vec_data_069_d2[1], vec_data_069_d2[2], vec_data_069_d2[3], vec_data_069_d2[4], vec_data_069_d2[5], vec_data_069_d2[6], vec_data_069_d2[7] };
  assign mask_d2_int16_w[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20905" *) { vec_data_070_d2[0], vec_data_070_d2[1], vec_data_070_d2[2], vec_data_070_d2[3], vec_data_070_d2[4], vec_data_070_d2[5], vec_data_070_d2[6], vec_data_070_d2[7], vec_data_071_d2[0], vec_data_071_d2[1], vec_data_071_d2[2], vec_data_071_d2[3], vec_data_071_d2[4], vec_data_071_d2[5], vec_data_071_d2[6], vec_data_071_d2[7] };
  assign mask_d2_int16_w[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20906" *) { vec_data_072_d2[0], vec_data_072_d2[1], vec_data_072_d2[2], vec_data_072_d2[3], vec_data_072_d2[4], vec_data_072_d2[5], vec_data_072_d2[6], vec_data_072_d2[7], vec_data_073_d2[0], vec_data_073_d2[1], vec_data_073_d2[2], vec_data_073_d2[3], vec_data_073_d2[4], vec_data_073_d2[5], vec_data_073_d2[6], vec_data_073_d2[7] };
  assign mask_d2_int16_w[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20907" *) { vec_data_074_d2[0], vec_data_074_d2[1], vec_data_074_d2[2], vec_data_074_d2[3], vec_data_074_d2[4], vec_data_074_d2[5], vec_data_074_d2[6], vec_data_074_d2[7], vec_data_075_d2[0], vec_data_075_d2[1], vec_data_075_d2[2], vec_data_075_d2[3], vec_data_075_d2[4], vec_data_075_d2[5], vec_data_075_d2[6], vec_data_075_d2[7] };
  assign mask_d2_int16_w[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20908" *) { vec_data_076_d2[0], vec_data_076_d2[1], vec_data_076_d2[2], vec_data_076_d2[3], vec_data_076_d2[4], vec_data_076_d2[5], vec_data_076_d2[6], vec_data_076_d2[7], vec_data_077_d2[0], vec_data_077_d2[1], vec_data_077_d2[2], vec_data_077_d2[3], vec_data_077_d2[4], vec_data_077_d2[5], vec_data_077_d2[6], vec_data_077_d2[7] };
  assign mask_d2_int16_w[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20909" *) { vec_data_078_d2[0], vec_data_078_d2[1], vec_data_078_d2[2], vec_data_078_d2[3], vec_data_078_d2[4], vec_data_078_d2[5], vec_data_078_d2[6], vec_data_078_d2[7], vec_data_079_d2[0], vec_data_079_d2[1], vec_data_079_d2[2], vec_data_079_d2[3], vec_data_079_d2[4], vec_data_079_d2[5], vec_data_079_d2[6], vec_data_079_d2[7] };
  assign mask_d2_int16_w[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20910" *) { vec_data_080_d2[0], vec_data_080_d2[1], vec_data_080_d2[2], vec_data_080_d2[3], vec_data_080_d2[4], vec_data_080_d2[5], vec_data_080_d2[6], vec_data_080_d2[7], vec_data_081_d2[0], vec_data_081_d2[1], vec_data_081_d2[2], vec_data_081_d2[3], vec_data_081_d2[4], vec_data_081_d2[5], vec_data_081_d2[6], vec_data_081_d2[7] };
  assign mask_d2_int16_w[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20911" *) { vec_data_082_d2[0], vec_data_082_d2[1], vec_data_082_d2[2], vec_data_082_d2[3], vec_data_082_d2[4], vec_data_082_d2[5], vec_data_082_d2[6], vec_data_082_d2[7], vec_data_083_d2[0], vec_data_083_d2[1], vec_data_083_d2[2], vec_data_083_d2[3], vec_data_083_d2[4], vec_data_083_d2[5], vec_data_083_d2[6], vec_data_083_d2[7] };
  assign mask_d2_int16_w[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20912" *) { vec_data_084_d2[0], vec_data_084_d2[1], vec_data_084_d2[2], vec_data_084_d2[3], vec_data_084_d2[4], vec_data_084_d2[5], vec_data_084_d2[6], vec_data_084_d2[7], vec_data_085_d2[0], vec_data_085_d2[1], vec_data_085_d2[2], vec_data_085_d2[3], vec_data_085_d2[4], vec_data_085_d2[5], vec_data_085_d2[6], vec_data_085_d2[7] };
  assign mask_d2_int16_w[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20913" *) { vec_data_086_d2[0], vec_data_086_d2[1], vec_data_086_d2[2], vec_data_086_d2[3], vec_data_086_d2[4], vec_data_086_d2[5], vec_data_086_d2[6], vec_data_086_d2[7], vec_data_087_d2[0], vec_data_087_d2[1], vec_data_087_d2[2], vec_data_087_d2[3], vec_data_087_d2[4], vec_data_087_d2[5], vec_data_087_d2[6], vec_data_087_d2[7] };
  assign mask_d2_int16_w[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20914" *) { vec_data_088_d2[0], vec_data_088_d2[1], vec_data_088_d2[2], vec_data_088_d2[3], vec_data_088_d2[4], vec_data_088_d2[5], vec_data_088_d2[6], vec_data_088_d2[7], vec_data_089_d2[0], vec_data_089_d2[1], vec_data_089_d2[2], vec_data_089_d2[3], vec_data_089_d2[4], vec_data_089_d2[5], vec_data_089_d2[6], vec_data_089_d2[7] };
  assign mask_d2_int16_w[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20915" *) { vec_data_090_d2[0], vec_data_090_d2[1], vec_data_090_d2[2], vec_data_090_d2[3], vec_data_090_d2[4], vec_data_090_d2[5], vec_data_090_d2[6], vec_data_090_d2[7], vec_data_091_d2[0], vec_data_091_d2[1], vec_data_091_d2[2], vec_data_091_d2[3], vec_data_091_d2[4], vec_data_091_d2[5], vec_data_091_d2[6], vec_data_091_d2[7] };
  assign mask_d2_int16_w[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20916" *) { vec_data_092_d2[0], vec_data_092_d2[1], vec_data_092_d2[2], vec_data_092_d2[3], vec_data_092_d2[4], vec_data_092_d2[5], vec_data_092_d2[6], vec_data_092_d2[7], vec_data_093_d2[0], vec_data_093_d2[1], vec_data_093_d2[2], vec_data_093_d2[3], vec_data_093_d2[4], vec_data_093_d2[5], vec_data_093_d2[6], vec_data_093_d2[7] };
  assign mask_d2_int16_w[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20917" *) { vec_data_094_d2[0], vec_data_094_d2[1], vec_data_094_d2[2], vec_data_094_d2[3], vec_data_094_d2[4], vec_data_094_d2[5], vec_data_094_d2[6], vec_data_094_d2[7], vec_data_095_d2[0], vec_data_095_d2[1], vec_data_095_d2[2], vec_data_095_d2[3], vec_data_095_d2[4], vec_data_095_d2[5], vec_data_095_d2[6], vec_data_095_d2[7] };
  assign mask_d2_int16_w[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20918" *) { vec_data_096_d2[0], vec_data_096_d2[1], vec_data_096_d2[2], vec_data_096_d2[3], vec_data_096_d2[4], vec_data_096_d2[5], vec_data_096_d2[6], vec_data_096_d2[7], vec_data_097_d2[0], vec_data_097_d2[1], vec_data_097_d2[2], vec_data_097_d2[3], vec_data_097_d2[4], vec_data_097_d2[5], vec_data_097_d2[6], vec_data_097_d2[7] };
  assign mask_d2_int16_w[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20919" *) { vec_data_098_d2[0], vec_data_098_d2[1], vec_data_098_d2[2], vec_data_098_d2[3], vec_data_098_d2[4], vec_data_098_d2[5], vec_data_098_d2[6], vec_data_098_d2[7], vec_data_099_d2[0], vec_data_099_d2[1], vec_data_099_d2[2], vec_data_099_d2[3], vec_data_099_d2[4], vec_data_099_d2[5], vec_data_099_d2[6], vec_data_099_d2[7] };
  assign mask_d2_int16_w[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20920" *) { vec_data_100_d2[0], vec_data_100_d2[1], vec_data_100_d2[2], vec_data_100_d2[3], vec_data_100_d2[4], vec_data_100_d2[5], vec_data_100_d2[6], vec_data_100_d2[7], vec_data_101_d2[0], vec_data_101_d2[1], vec_data_101_d2[2], vec_data_101_d2[3], vec_data_101_d2[4], vec_data_101_d2[5], vec_data_101_d2[6], vec_data_101_d2[7] };
  assign mask_d2_int16_w[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20921" *) { vec_data_102_d2[0], vec_data_102_d2[1], vec_data_102_d2[2], vec_data_102_d2[3], vec_data_102_d2[4], vec_data_102_d2[5], vec_data_102_d2[6], vec_data_102_d2[7], vec_data_103_d2[0], vec_data_103_d2[1], vec_data_103_d2[2], vec_data_103_d2[3], vec_data_103_d2[4], vec_data_103_d2[5], vec_data_103_d2[6], vec_data_103_d2[7] };
  assign mask_d2_int16_w[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20922" *) { vec_data_104_d2[0], vec_data_104_d2[1], vec_data_104_d2[2], vec_data_104_d2[3], vec_data_104_d2[4], vec_data_104_d2[5], vec_data_104_d2[6], vec_data_104_d2[7], vec_data_105_d2[0], vec_data_105_d2[1], vec_data_105_d2[2], vec_data_105_d2[3], vec_data_105_d2[4], vec_data_105_d2[5], vec_data_105_d2[6], vec_data_105_d2[7] };
  assign mask_d2_int16_w[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20923" *) { vec_data_106_d2[0], vec_data_106_d2[1], vec_data_106_d2[2], vec_data_106_d2[3], vec_data_106_d2[4], vec_data_106_d2[5], vec_data_106_d2[6], vec_data_106_d2[7], vec_data_107_d2[0], vec_data_107_d2[1], vec_data_107_d2[2], vec_data_107_d2[3], vec_data_107_d2[4], vec_data_107_d2[5], vec_data_107_d2[6], vec_data_107_d2[7] };
  assign mask_d2_int16_w[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20924" *) { vec_data_108_d2[0], vec_data_108_d2[1], vec_data_108_d2[2], vec_data_108_d2[3], vec_data_108_d2[4], vec_data_108_d2[5], vec_data_108_d2[6], vec_data_108_d2[7], vec_data_109_d2[0], vec_data_109_d2[1], vec_data_109_d2[2], vec_data_109_d2[3], vec_data_109_d2[4], vec_data_109_d2[5], vec_data_109_d2[6], vec_data_109_d2[7] };
  assign mask_d2_int16_w[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20925" *) { vec_data_110_d2[0], vec_data_110_d2[1], vec_data_110_d2[2], vec_data_110_d2[3], vec_data_110_d2[4], vec_data_110_d2[5], vec_data_110_d2[6], vec_data_110_d2[7], vec_data_111_d2[0], vec_data_111_d2[1], vec_data_111_d2[2], vec_data_111_d2[3], vec_data_111_d2[4], vec_data_111_d2[5], vec_data_111_d2[6], vec_data_111_d2[7] };
  assign mask_d2_int16_w[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20926" *) { vec_data_112_d2[0], vec_data_112_d2[1], vec_data_112_d2[2], vec_data_112_d2[3], vec_data_112_d2[4], vec_data_112_d2[5], vec_data_112_d2[6], vec_data_112_d2[7], vec_data_113_d2[0], vec_data_113_d2[1], vec_data_113_d2[2], vec_data_113_d2[3], vec_data_113_d2[4], vec_data_113_d2[5], vec_data_113_d2[6], vec_data_113_d2[7] };
  assign mask_d2_int16_w[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20927" *) { vec_data_114_d2[0], vec_data_114_d2[1], vec_data_114_d2[2], vec_data_114_d2[3], vec_data_114_d2[4], vec_data_114_d2[5], vec_data_114_d2[6], vec_data_114_d2[7], vec_data_115_d2[0], vec_data_115_d2[1], vec_data_115_d2[2], vec_data_115_d2[3], vec_data_115_d2[4], vec_data_115_d2[5], vec_data_115_d2[6], vec_data_115_d2[7] };
  assign mask_d2_int16_w[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20928" *) { vec_data_116_d2[0], vec_data_116_d2[1], vec_data_116_d2[2], vec_data_116_d2[3], vec_data_116_d2[4], vec_data_116_d2[5], vec_data_116_d2[6], vec_data_116_d2[7], vec_data_117_d2[0], vec_data_117_d2[1], vec_data_117_d2[2], vec_data_117_d2[3], vec_data_117_d2[4], vec_data_117_d2[5], vec_data_117_d2[6], vec_data_117_d2[7] };
  assign mask_d2_int16_w[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20929" *) { vec_data_118_d2[0], vec_data_118_d2[1], vec_data_118_d2[2], vec_data_118_d2[3], vec_data_118_d2[4], vec_data_118_d2[5], vec_data_118_d2[6], vec_data_118_d2[7], vec_data_119_d2[0], vec_data_119_d2[1], vec_data_119_d2[2], vec_data_119_d2[3], vec_data_119_d2[4], vec_data_119_d2[5], vec_data_119_d2[6], vec_data_119_d2[7] };
  assign mask_d2_int16_w[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20930" *) { vec_data_120_d2[0], vec_data_120_d2[1], vec_data_120_d2[2], vec_data_120_d2[3], vec_data_120_d2[4], vec_data_120_d2[5], vec_data_120_d2[6], vec_data_120_d2[7], vec_data_121_d2[0], vec_data_121_d2[1], vec_data_121_d2[2], vec_data_121_d2[3], vec_data_121_d2[4], vec_data_121_d2[5], vec_data_121_d2[6], vec_data_121_d2[7] };
  assign mask_d2_int16_w[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20931" *) { vec_data_122_d2[0], vec_data_122_d2[1], vec_data_122_d2[2], vec_data_122_d2[3], vec_data_122_d2[4], vec_data_122_d2[5], vec_data_122_d2[6], vec_data_122_d2[7], vec_data_123_d2[0], vec_data_123_d2[1], vec_data_123_d2[2], vec_data_123_d2[3], vec_data_123_d2[4], vec_data_123_d2[5], vec_data_123_d2[6], vec_data_123_d2[7] };
  assign mask_d2_int16_w[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20932" *) { vec_data_124_d2[0], vec_data_124_d2[1], vec_data_124_d2[2], vec_data_124_d2[3], vec_data_124_d2[4], vec_data_124_d2[5], vec_data_124_d2[6], vec_data_124_d2[7], vec_data_125_d2[0], vec_data_125_d2[1], vec_data_125_d2[2], vec_data_125_d2[3], vec_data_125_d2[4], vec_data_125_d2[5], vec_data_125_d2[6], vec_data_125_d2[7] };
  assign mask_d2_int16_w[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:20933" *) { vec_data_126_d2[0], vec_data_126_d2[1], vec_data_126_d2[2], vec_data_126_d2[3], vec_data_126_d2[4], vec_data_126_d2[5], vec_data_126_d2[6], vec_data_126_d2[7], vec_data_127_d2[0], vec_data_127_d2[1], vec_data_127_d2[2], vec_data_127_d2[3], vec_data_127_d2[4], vec_data_127_d2[5], vec_data_127_d2[6], vec_data_127_d2[7] };
  assign mask_d2_fp16_w[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21065" *) { vec_data_000_d2[0], vec_data_000_d2[1], vec_data_000_d2[2], vec_data_000_d2[3], vec_data_000_d2[4], vec_data_000_d2[5], vec_data_000_d2[6], vec_data_000_d2[7], vec_data_001_d2[0], vec_data_001_d2[1], vec_data_001_d2[2], vec_data_001_d2[3], vec_data_001_d2[4], vec_data_001_d2[5], vec_data_001_d2[6] };
  assign mask_d2_fp16_w[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21066" *) { vec_data_002_d2[0], vec_data_002_d2[1], vec_data_002_d2[2], vec_data_002_d2[3], vec_data_002_d2[4], vec_data_002_d2[5], vec_data_002_d2[6], vec_data_002_d2[7], vec_data_003_d2[0], vec_data_003_d2[1], vec_data_003_d2[2], vec_data_003_d2[3], vec_data_003_d2[4], vec_data_003_d2[5], vec_data_003_d2[6] };
  assign mask_d2_fp16_w[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21067" *) { vec_data_004_d2[0], vec_data_004_d2[1], vec_data_004_d2[2], vec_data_004_d2[3], vec_data_004_d2[4], vec_data_004_d2[5], vec_data_004_d2[6], vec_data_004_d2[7], vec_data_005_d2[0], vec_data_005_d2[1], vec_data_005_d2[2], vec_data_005_d2[3], vec_data_005_d2[4], vec_data_005_d2[5], vec_data_005_d2[6] };
  assign mask_d2_fp16_w[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21068" *) { vec_data_006_d2[0], vec_data_006_d2[1], vec_data_006_d2[2], vec_data_006_d2[3], vec_data_006_d2[4], vec_data_006_d2[5], vec_data_006_d2[6], vec_data_006_d2[7], vec_data_007_d2[0], vec_data_007_d2[1], vec_data_007_d2[2], vec_data_007_d2[3], vec_data_007_d2[4], vec_data_007_d2[5], vec_data_007_d2[6] };
  assign mask_d2_fp16_w[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21069" *) { vec_data_008_d2[0], vec_data_008_d2[1], vec_data_008_d2[2], vec_data_008_d2[3], vec_data_008_d2[4], vec_data_008_d2[5], vec_data_008_d2[6], vec_data_008_d2[7], vec_data_009_d2[0], vec_data_009_d2[1], vec_data_009_d2[2], vec_data_009_d2[3], vec_data_009_d2[4], vec_data_009_d2[5], vec_data_009_d2[6] };
  assign mask_d2_fp16_w[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21070" *) { vec_data_010_d2[0], vec_data_010_d2[1], vec_data_010_d2[2], vec_data_010_d2[3], vec_data_010_d2[4], vec_data_010_d2[5], vec_data_010_d2[6], vec_data_010_d2[7], vec_data_011_d2[0], vec_data_011_d2[1], vec_data_011_d2[2], vec_data_011_d2[3], vec_data_011_d2[4], vec_data_011_d2[5], vec_data_011_d2[6] };
  assign mask_d2_fp16_w[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21071" *) { vec_data_012_d2[0], vec_data_012_d2[1], vec_data_012_d2[2], vec_data_012_d2[3], vec_data_012_d2[4], vec_data_012_d2[5], vec_data_012_d2[6], vec_data_012_d2[7], vec_data_013_d2[0], vec_data_013_d2[1], vec_data_013_d2[2], vec_data_013_d2[3], vec_data_013_d2[4], vec_data_013_d2[5], vec_data_013_d2[6] };
  assign mask_d2_fp16_w[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21072" *) { vec_data_014_d2[0], vec_data_014_d2[1], vec_data_014_d2[2], vec_data_014_d2[3], vec_data_014_d2[4], vec_data_014_d2[5], vec_data_014_d2[6], vec_data_014_d2[7], vec_data_015_d2[0], vec_data_015_d2[1], vec_data_015_d2[2], vec_data_015_d2[3], vec_data_015_d2[4], vec_data_015_d2[5], vec_data_015_d2[6] };
  assign mask_d2_fp16_w[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21073" *) { vec_data_016_d2[0], vec_data_016_d2[1], vec_data_016_d2[2], vec_data_016_d2[3], vec_data_016_d2[4], vec_data_016_d2[5], vec_data_016_d2[6], vec_data_016_d2[7], vec_data_017_d2[0], vec_data_017_d2[1], vec_data_017_d2[2], vec_data_017_d2[3], vec_data_017_d2[4], vec_data_017_d2[5], vec_data_017_d2[6] };
  assign mask_d2_fp16_w[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21074" *) { vec_data_018_d2[0], vec_data_018_d2[1], vec_data_018_d2[2], vec_data_018_d2[3], vec_data_018_d2[4], vec_data_018_d2[5], vec_data_018_d2[6], vec_data_018_d2[7], vec_data_019_d2[0], vec_data_019_d2[1], vec_data_019_d2[2], vec_data_019_d2[3], vec_data_019_d2[4], vec_data_019_d2[5], vec_data_019_d2[6] };
  assign mask_d2_fp16_w[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21075" *) { vec_data_020_d2[0], vec_data_020_d2[1], vec_data_020_d2[2], vec_data_020_d2[3], vec_data_020_d2[4], vec_data_020_d2[5], vec_data_020_d2[6], vec_data_020_d2[7], vec_data_021_d2[0], vec_data_021_d2[1], vec_data_021_d2[2], vec_data_021_d2[3], vec_data_021_d2[4], vec_data_021_d2[5], vec_data_021_d2[6] };
  assign mask_d2_fp16_w[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21076" *) { vec_data_022_d2[0], vec_data_022_d2[1], vec_data_022_d2[2], vec_data_022_d2[3], vec_data_022_d2[4], vec_data_022_d2[5], vec_data_022_d2[6], vec_data_022_d2[7], vec_data_023_d2[0], vec_data_023_d2[1], vec_data_023_d2[2], vec_data_023_d2[3], vec_data_023_d2[4], vec_data_023_d2[5], vec_data_023_d2[6] };
  assign mask_d2_fp16_w[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21077" *) { vec_data_024_d2[0], vec_data_024_d2[1], vec_data_024_d2[2], vec_data_024_d2[3], vec_data_024_d2[4], vec_data_024_d2[5], vec_data_024_d2[6], vec_data_024_d2[7], vec_data_025_d2[0], vec_data_025_d2[1], vec_data_025_d2[2], vec_data_025_d2[3], vec_data_025_d2[4], vec_data_025_d2[5], vec_data_025_d2[6] };
  assign mask_d2_fp16_w[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21078" *) { vec_data_026_d2[0], vec_data_026_d2[1], vec_data_026_d2[2], vec_data_026_d2[3], vec_data_026_d2[4], vec_data_026_d2[5], vec_data_026_d2[6], vec_data_026_d2[7], vec_data_027_d2[0], vec_data_027_d2[1], vec_data_027_d2[2], vec_data_027_d2[3], vec_data_027_d2[4], vec_data_027_d2[5], vec_data_027_d2[6] };
  assign mask_d2_fp16_w[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21079" *) { vec_data_028_d2[0], vec_data_028_d2[1], vec_data_028_d2[2], vec_data_028_d2[3], vec_data_028_d2[4], vec_data_028_d2[5], vec_data_028_d2[6], vec_data_028_d2[7], vec_data_029_d2[0], vec_data_029_d2[1], vec_data_029_d2[2], vec_data_029_d2[3], vec_data_029_d2[4], vec_data_029_d2[5], vec_data_029_d2[6] };
  assign mask_d2_fp16_w[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21080" *) { vec_data_030_d2[0], vec_data_030_d2[1], vec_data_030_d2[2], vec_data_030_d2[3], vec_data_030_d2[4], vec_data_030_d2[5], vec_data_030_d2[6], vec_data_030_d2[7], vec_data_031_d2[0], vec_data_031_d2[1], vec_data_031_d2[2], vec_data_031_d2[3], vec_data_031_d2[4], vec_data_031_d2[5], vec_data_031_d2[6] };
  assign mask_d2_fp16_w[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21081" *) { vec_data_032_d2[0], vec_data_032_d2[1], vec_data_032_d2[2], vec_data_032_d2[3], vec_data_032_d2[4], vec_data_032_d2[5], vec_data_032_d2[6], vec_data_032_d2[7], vec_data_033_d2[0], vec_data_033_d2[1], vec_data_033_d2[2], vec_data_033_d2[3], vec_data_033_d2[4], vec_data_033_d2[5], vec_data_033_d2[6] };
  assign mask_d2_fp16_w[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21082" *) { vec_data_034_d2[0], vec_data_034_d2[1], vec_data_034_d2[2], vec_data_034_d2[3], vec_data_034_d2[4], vec_data_034_d2[5], vec_data_034_d2[6], vec_data_034_d2[7], vec_data_035_d2[0], vec_data_035_d2[1], vec_data_035_d2[2], vec_data_035_d2[3], vec_data_035_d2[4], vec_data_035_d2[5], vec_data_035_d2[6] };
  assign mask_d2_fp16_w[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21083" *) { vec_data_036_d2[0], vec_data_036_d2[1], vec_data_036_d2[2], vec_data_036_d2[3], vec_data_036_d2[4], vec_data_036_d2[5], vec_data_036_d2[6], vec_data_036_d2[7], vec_data_037_d2[0], vec_data_037_d2[1], vec_data_037_d2[2], vec_data_037_d2[3], vec_data_037_d2[4], vec_data_037_d2[5], vec_data_037_d2[6] };
  assign mask_d2_fp16_w[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21084" *) { vec_data_038_d2[0], vec_data_038_d2[1], vec_data_038_d2[2], vec_data_038_d2[3], vec_data_038_d2[4], vec_data_038_d2[5], vec_data_038_d2[6], vec_data_038_d2[7], vec_data_039_d2[0], vec_data_039_d2[1], vec_data_039_d2[2], vec_data_039_d2[3], vec_data_039_d2[4], vec_data_039_d2[5], vec_data_039_d2[6] };
  assign mask_d2_fp16_w[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21085" *) { vec_data_040_d2[0], vec_data_040_d2[1], vec_data_040_d2[2], vec_data_040_d2[3], vec_data_040_d2[4], vec_data_040_d2[5], vec_data_040_d2[6], vec_data_040_d2[7], vec_data_041_d2[0], vec_data_041_d2[1], vec_data_041_d2[2], vec_data_041_d2[3], vec_data_041_d2[4], vec_data_041_d2[5], vec_data_041_d2[6] };
  assign mask_d2_fp16_w[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21086" *) { vec_data_042_d2[0], vec_data_042_d2[1], vec_data_042_d2[2], vec_data_042_d2[3], vec_data_042_d2[4], vec_data_042_d2[5], vec_data_042_d2[6], vec_data_042_d2[7], vec_data_043_d2[0], vec_data_043_d2[1], vec_data_043_d2[2], vec_data_043_d2[3], vec_data_043_d2[4], vec_data_043_d2[5], vec_data_043_d2[6] };
  assign mask_d2_fp16_w[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21087" *) { vec_data_044_d2[0], vec_data_044_d2[1], vec_data_044_d2[2], vec_data_044_d2[3], vec_data_044_d2[4], vec_data_044_d2[5], vec_data_044_d2[6], vec_data_044_d2[7], vec_data_045_d2[0], vec_data_045_d2[1], vec_data_045_d2[2], vec_data_045_d2[3], vec_data_045_d2[4], vec_data_045_d2[5], vec_data_045_d2[6] };
  assign mask_d2_fp16_w[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21088" *) { vec_data_046_d2[0], vec_data_046_d2[1], vec_data_046_d2[2], vec_data_046_d2[3], vec_data_046_d2[4], vec_data_046_d2[5], vec_data_046_d2[6], vec_data_046_d2[7], vec_data_047_d2[0], vec_data_047_d2[1], vec_data_047_d2[2], vec_data_047_d2[3], vec_data_047_d2[4], vec_data_047_d2[5], vec_data_047_d2[6] };
  assign mask_d2_fp16_w[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21089" *) { vec_data_048_d2[0], vec_data_048_d2[1], vec_data_048_d2[2], vec_data_048_d2[3], vec_data_048_d2[4], vec_data_048_d2[5], vec_data_048_d2[6], vec_data_048_d2[7], vec_data_049_d2[0], vec_data_049_d2[1], vec_data_049_d2[2], vec_data_049_d2[3], vec_data_049_d2[4], vec_data_049_d2[5], vec_data_049_d2[6] };
  assign mask_d2_fp16_w[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21090" *) { vec_data_050_d2[0], vec_data_050_d2[1], vec_data_050_d2[2], vec_data_050_d2[3], vec_data_050_d2[4], vec_data_050_d2[5], vec_data_050_d2[6], vec_data_050_d2[7], vec_data_051_d2[0], vec_data_051_d2[1], vec_data_051_d2[2], vec_data_051_d2[3], vec_data_051_d2[4], vec_data_051_d2[5], vec_data_051_d2[6] };
  assign mask_d2_fp16_w[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21091" *) { vec_data_052_d2[0], vec_data_052_d2[1], vec_data_052_d2[2], vec_data_052_d2[3], vec_data_052_d2[4], vec_data_052_d2[5], vec_data_052_d2[6], vec_data_052_d2[7], vec_data_053_d2[0], vec_data_053_d2[1], vec_data_053_d2[2], vec_data_053_d2[3], vec_data_053_d2[4], vec_data_053_d2[5], vec_data_053_d2[6] };
  assign mask_d2_fp16_w[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21092" *) { vec_data_054_d2[0], vec_data_054_d2[1], vec_data_054_d2[2], vec_data_054_d2[3], vec_data_054_d2[4], vec_data_054_d2[5], vec_data_054_d2[6], vec_data_054_d2[7], vec_data_055_d2[0], vec_data_055_d2[1], vec_data_055_d2[2], vec_data_055_d2[3], vec_data_055_d2[4], vec_data_055_d2[5], vec_data_055_d2[6] };
  assign mask_d2_fp16_w[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21093" *) { vec_data_056_d2[0], vec_data_056_d2[1], vec_data_056_d2[2], vec_data_056_d2[3], vec_data_056_d2[4], vec_data_056_d2[5], vec_data_056_d2[6], vec_data_056_d2[7], vec_data_057_d2[0], vec_data_057_d2[1], vec_data_057_d2[2], vec_data_057_d2[3], vec_data_057_d2[4], vec_data_057_d2[5], vec_data_057_d2[6] };
  assign mask_d2_fp16_w[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21094" *) { vec_data_058_d2[0], vec_data_058_d2[1], vec_data_058_d2[2], vec_data_058_d2[3], vec_data_058_d2[4], vec_data_058_d2[5], vec_data_058_d2[6], vec_data_058_d2[7], vec_data_059_d2[0], vec_data_059_d2[1], vec_data_059_d2[2], vec_data_059_d2[3], vec_data_059_d2[4], vec_data_059_d2[5], vec_data_059_d2[6] };
  assign mask_d2_fp16_w[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21095" *) { vec_data_060_d2[0], vec_data_060_d2[1], vec_data_060_d2[2], vec_data_060_d2[3], vec_data_060_d2[4], vec_data_060_d2[5], vec_data_060_d2[6], vec_data_060_d2[7], vec_data_061_d2[0], vec_data_061_d2[1], vec_data_061_d2[2], vec_data_061_d2[3], vec_data_061_d2[4], vec_data_061_d2[5], vec_data_061_d2[6] };
  assign mask_d2_fp16_w[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21096" *) { vec_data_062_d2[0], vec_data_062_d2[1], vec_data_062_d2[2], vec_data_062_d2[3], vec_data_062_d2[4], vec_data_062_d2[5], vec_data_062_d2[6], vec_data_062_d2[7], vec_data_063_d2[0], vec_data_063_d2[1], vec_data_063_d2[2], vec_data_063_d2[3], vec_data_063_d2[4], vec_data_063_d2[5], vec_data_063_d2[6] };
  assign mask_d2_fp16_w[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21097" *) { vec_data_064_d2[0], vec_data_064_d2[1], vec_data_064_d2[2], vec_data_064_d2[3], vec_data_064_d2[4], vec_data_064_d2[5], vec_data_064_d2[6], vec_data_064_d2[7], vec_data_065_d2[0], vec_data_065_d2[1], vec_data_065_d2[2], vec_data_065_d2[3], vec_data_065_d2[4], vec_data_065_d2[5], vec_data_065_d2[6] };
  assign mask_d2_fp16_w[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21098" *) { vec_data_066_d2[0], vec_data_066_d2[1], vec_data_066_d2[2], vec_data_066_d2[3], vec_data_066_d2[4], vec_data_066_d2[5], vec_data_066_d2[6], vec_data_066_d2[7], vec_data_067_d2[0], vec_data_067_d2[1], vec_data_067_d2[2], vec_data_067_d2[3], vec_data_067_d2[4], vec_data_067_d2[5], vec_data_067_d2[6] };
  assign mask_d2_fp16_w[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21099" *) { vec_data_068_d2[0], vec_data_068_d2[1], vec_data_068_d2[2], vec_data_068_d2[3], vec_data_068_d2[4], vec_data_068_d2[5], vec_data_068_d2[6], vec_data_068_d2[7], vec_data_069_d2[0], vec_data_069_d2[1], vec_data_069_d2[2], vec_data_069_d2[3], vec_data_069_d2[4], vec_data_069_d2[5], vec_data_069_d2[6] };
  assign mask_d2_fp16_w[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21100" *) { vec_data_070_d2[0], vec_data_070_d2[1], vec_data_070_d2[2], vec_data_070_d2[3], vec_data_070_d2[4], vec_data_070_d2[5], vec_data_070_d2[6], vec_data_070_d2[7], vec_data_071_d2[0], vec_data_071_d2[1], vec_data_071_d2[2], vec_data_071_d2[3], vec_data_071_d2[4], vec_data_071_d2[5], vec_data_071_d2[6] };
  assign mask_d2_fp16_w[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21101" *) { vec_data_072_d2[0], vec_data_072_d2[1], vec_data_072_d2[2], vec_data_072_d2[3], vec_data_072_d2[4], vec_data_072_d2[5], vec_data_072_d2[6], vec_data_072_d2[7], vec_data_073_d2[0], vec_data_073_d2[1], vec_data_073_d2[2], vec_data_073_d2[3], vec_data_073_d2[4], vec_data_073_d2[5], vec_data_073_d2[6] };
  assign mask_d2_fp16_w[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21102" *) { vec_data_074_d2[0], vec_data_074_d2[1], vec_data_074_d2[2], vec_data_074_d2[3], vec_data_074_d2[4], vec_data_074_d2[5], vec_data_074_d2[6], vec_data_074_d2[7], vec_data_075_d2[0], vec_data_075_d2[1], vec_data_075_d2[2], vec_data_075_d2[3], vec_data_075_d2[4], vec_data_075_d2[5], vec_data_075_d2[6] };
  assign mask_d2_fp16_w[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21103" *) { vec_data_076_d2[0], vec_data_076_d2[1], vec_data_076_d2[2], vec_data_076_d2[3], vec_data_076_d2[4], vec_data_076_d2[5], vec_data_076_d2[6], vec_data_076_d2[7], vec_data_077_d2[0], vec_data_077_d2[1], vec_data_077_d2[2], vec_data_077_d2[3], vec_data_077_d2[4], vec_data_077_d2[5], vec_data_077_d2[6] };
  assign mask_d2_fp16_w[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21104" *) { vec_data_078_d2[0], vec_data_078_d2[1], vec_data_078_d2[2], vec_data_078_d2[3], vec_data_078_d2[4], vec_data_078_d2[5], vec_data_078_d2[6], vec_data_078_d2[7], vec_data_079_d2[0], vec_data_079_d2[1], vec_data_079_d2[2], vec_data_079_d2[3], vec_data_079_d2[4], vec_data_079_d2[5], vec_data_079_d2[6] };
  assign mask_d2_fp16_w[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21105" *) { vec_data_080_d2[0], vec_data_080_d2[1], vec_data_080_d2[2], vec_data_080_d2[3], vec_data_080_d2[4], vec_data_080_d2[5], vec_data_080_d2[6], vec_data_080_d2[7], vec_data_081_d2[0], vec_data_081_d2[1], vec_data_081_d2[2], vec_data_081_d2[3], vec_data_081_d2[4], vec_data_081_d2[5], vec_data_081_d2[6] };
  assign mask_d2_fp16_w[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21106" *) { vec_data_082_d2[0], vec_data_082_d2[1], vec_data_082_d2[2], vec_data_082_d2[3], vec_data_082_d2[4], vec_data_082_d2[5], vec_data_082_d2[6], vec_data_082_d2[7], vec_data_083_d2[0], vec_data_083_d2[1], vec_data_083_d2[2], vec_data_083_d2[3], vec_data_083_d2[4], vec_data_083_d2[5], vec_data_083_d2[6] };
  assign mask_d2_fp16_w[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21107" *) { vec_data_084_d2[0], vec_data_084_d2[1], vec_data_084_d2[2], vec_data_084_d2[3], vec_data_084_d2[4], vec_data_084_d2[5], vec_data_084_d2[6], vec_data_084_d2[7], vec_data_085_d2[0], vec_data_085_d2[1], vec_data_085_d2[2], vec_data_085_d2[3], vec_data_085_d2[4], vec_data_085_d2[5], vec_data_085_d2[6] };
  assign mask_d2_fp16_w[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21108" *) { vec_data_086_d2[0], vec_data_086_d2[1], vec_data_086_d2[2], vec_data_086_d2[3], vec_data_086_d2[4], vec_data_086_d2[5], vec_data_086_d2[6], vec_data_086_d2[7], vec_data_087_d2[0], vec_data_087_d2[1], vec_data_087_d2[2], vec_data_087_d2[3], vec_data_087_d2[4], vec_data_087_d2[5], vec_data_087_d2[6] };
  assign mask_d2_fp16_w[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21109" *) { vec_data_088_d2[0], vec_data_088_d2[1], vec_data_088_d2[2], vec_data_088_d2[3], vec_data_088_d2[4], vec_data_088_d2[5], vec_data_088_d2[6], vec_data_088_d2[7], vec_data_089_d2[0], vec_data_089_d2[1], vec_data_089_d2[2], vec_data_089_d2[3], vec_data_089_d2[4], vec_data_089_d2[5], vec_data_089_d2[6] };
  assign mask_d2_fp16_w[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21110" *) { vec_data_090_d2[0], vec_data_090_d2[1], vec_data_090_d2[2], vec_data_090_d2[3], vec_data_090_d2[4], vec_data_090_d2[5], vec_data_090_d2[6], vec_data_090_d2[7], vec_data_091_d2[0], vec_data_091_d2[1], vec_data_091_d2[2], vec_data_091_d2[3], vec_data_091_d2[4], vec_data_091_d2[5], vec_data_091_d2[6] };
  assign mask_d2_fp16_w[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21111" *) { vec_data_092_d2[0], vec_data_092_d2[1], vec_data_092_d2[2], vec_data_092_d2[3], vec_data_092_d2[4], vec_data_092_d2[5], vec_data_092_d2[6], vec_data_092_d2[7], vec_data_093_d2[0], vec_data_093_d2[1], vec_data_093_d2[2], vec_data_093_d2[3], vec_data_093_d2[4], vec_data_093_d2[5], vec_data_093_d2[6] };
  assign mask_d2_fp16_w[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21112" *) { vec_data_094_d2[0], vec_data_094_d2[1], vec_data_094_d2[2], vec_data_094_d2[3], vec_data_094_d2[4], vec_data_094_d2[5], vec_data_094_d2[6], vec_data_094_d2[7], vec_data_095_d2[0], vec_data_095_d2[1], vec_data_095_d2[2], vec_data_095_d2[3], vec_data_095_d2[4], vec_data_095_d2[5], vec_data_095_d2[6] };
  assign mask_d2_fp16_w[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21113" *) { vec_data_096_d2[0], vec_data_096_d2[1], vec_data_096_d2[2], vec_data_096_d2[3], vec_data_096_d2[4], vec_data_096_d2[5], vec_data_096_d2[6], vec_data_096_d2[7], vec_data_097_d2[0], vec_data_097_d2[1], vec_data_097_d2[2], vec_data_097_d2[3], vec_data_097_d2[4], vec_data_097_d2[5], vec_data_097_d2[6] };
  assign mask_d2_fp16_w[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21114" *) { vec_data_098_d2[0], vec_data_098_d2[1], vec_data_098_d2[2], vec_data_098_d2[3], vec_data_098_d2[4], vec_data_098_d2[5], vec_data_098_d2[6], vec_data_098_d2[7], vec_data_099_d2[0], vec_data_099_d2[1], vec_data_099_d2[2], vec_data_099_d2[3], vec_data_099_d2[4], vec_data_099_d2[5], vec_data_099_d2[6] };
  assign mask_d2_fp16_w[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21115" *) { vec_data_100_d2[0], vec_data_100_d2[1], vec_data_100_d2[2], vec_data_100_d2[3], vec_data_100_d2[4], vec_data_100_d2[5], vec_data_100_d2[6], vec_data_100_d2[7], vec_data_101_d2[0], vec_data_101_d2[1], vec_data_101_d2[2], vec_data_101_d2[3], vec_data_101_d2[4], vec_data_101_d2[5], vec_data_101_d2[6] };
  assign mask_d2_fp16_w[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21116" *) { vec_data_102_d2[0], vec_data_102_d2[1], vec_data_102_d2[2], vec_data_102_d2[3], vec_data_102_d2[4], vec_data_102_d2[5], vec_data_102_d2[6], vec_data_102_d2[7], vec_data_103_d2[0], vec_data_103_d2[1], vec_data_103_d2[2], vec_data_103_d2[3], vec_data_103_d2[4], vec_data_103_d2[5], vec_data_103_d2[6] };
  assign mask_d2_fp16_w[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21117" *) { vec_data_104_d2[0], vec_data_104_d2[1], vec_data_104_d2[2], vec_data_104_d2[3], vec_data_104_d2[4], vec_data_104_d2[5], vec_data_104_d2[6], vec_data_104_d2[7], vec_data_105_d2[0], vec_data_105_d2[1], vec_data_105_d2[2], vec_data_105_d2[3], vec_data_105_d2[4], vec_data_105_d2[5], vec_data_105_d2[6] };
  assign mask_d2_fp16_w[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21118" *) { vec_data_106_d2[0], vec_data_106_d2[1], vec_data_106_d2[2], vec_data_106_d2[3], vec_data_106_d2[4], vec_data_106_d2[5], vec_data_106_d2[6], vec_data_106_d2[7], vec_data_107_d2[0], vec_data_107_d2[1], vec_data_107_d2[2], vec_data_107_d2[3], vec_data_107_d2[4], vec_data_107_d2[5], vec_data_107_d2[6] };
  assign mask_d2_fp16_w[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21119" *) { vec_data_108_d2[0], vec_data_108_d2[1], vec_data_108_d2[2], vec_data_108_d2[3], vec_data_108_d2[4], vec_data_108_d2[5], vec_data_108_d2[6], vec_data_108_d2[7], vec_data_109_d2[0], vec_data_109_d2[1], vec_data_109_d2[2], vec_data_109_d2[3], vec_data_109_d2[4], vec_data_109_d2[5], vec_data_109_d2[6] };
  assign mask_d2_fp16_w[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21120" *) { vec_data_110_d2[0], vec_data_110_d2[1], vec_data_110_d2[2], vec_data_110_d2[3], vec_data_110_d2[4], vec_data_110_d2[5], vec_data_110_d2[6], vec_data_110_d2[7], vec_data_111_d2[0], vec_data_111_d2[1], vec_data_111_d2[2], vec_data_111_d2[3], vec_data_111_d2[4], vec_data_111_d2[5], vec_data_111_d2[6] };
  assign mask_d2_fp16_w[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21121" *) { vec_data_112_d2[0], vec_data_112_d2[1], vec_data_112_d2[2], vec_data_112_d2[3], vec_data_112_d2[4], vec_data_112_d2[5], vec_data_112_d2[6], vec_data_112_d2[7], vec_data_113_d2[0], vec_data_113_d2[1], vec_data_113_d2[2], vec_data_113_d2[3], vec_data_113_d2[4], vec_data_113_d2[5], vec_data_113_d2[6] };
  assign mask_d2_fp16_w[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21122" *) { vec_data_114_d2[0], vec_data_114_d2[1], vec_data_114_d2[2], vec_data_114_d2[3], vec_data_114_d2[4], vec_data_114_d2[5], vec_data_114_d2[6], vec_data_114_d2[7], vec_data_115_d2[0], vec_data_115_d2[1], vec_data_115_d2[2], vec_data_115_d2[3], vec_data_115_d2[4], vec_data_115_d2[5], vec_data_115_d2[6] };
  assign mask_d2_fp16_w[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21123" *) { vec_data_116_d2[0], vec_data_116_d2[1], vec_data_116_d2[2], vec_data_116_d2[3], vec_data_116_d2[4], vec_data_116_d2[5], vec_data_116_d2[6], vec_data_116_d2[7], vec_data_117_d2[0], vec_data_117_d2[1], vec_data_117_d2[2], vec_data_117_d2[3], vec_data_117_d2[4], vec_data_117_d2[5], vec_data_117_d2[6] };
  assign mask_d2_fp16_w[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21124" *) { vec_data_118_d2[0], vec_data_118_d2[1], vec_data_118_d2[2], vec_data_118_d2[3], vec_data_118_d2[4], vec_data_118_d2[5], vec_data_118_d2[6], vec_data_118_d2[7], vec_data_119_d2[0], vec_data_119_d2[1], vec_data_119_d2[2], vec_data_119_d2[3], vec_data_119_d2[4], vec_data_119_d2[5], vec_data_119_d2[6] };
  assign mask_d2_fp16_w[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21125" *) { vec_data_120_d2[0], vec_data_120_d2[1], vec_data_120_d2[2], vec_data_120_d2[3], vec_data_120_d2[4], vec_data_120_d2[5], vec_data_120_d2[6], vec_data_120_d2[7], vec_data_121_d2[0], vec_data_121_d2[1], vec_data_121_d2[2], vec_data_121_d2[3], vec_data_121_d2[4], vec_data_121_d2[5], vec_data_121_d2[6] };
  assign mask_d2_fp16_w[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21126" *) { vec_data_122_d2[0], vec_data_122_d2[1], vec_data_122_d2[2], vec_data_122_d2[3], vec_data_122_d2[4], vec_data_122_d2[5], vec_data_122_d2[6], vec_data_122_d2[7], vec_data_123_d2[0], vec_data_123_d2[1], vec_data_123_d2[2], vec_data_123_d2[3], vec_data_123_d2[4], vec_data_123_d2[5], vec_data_123_d2[6] };
  assign mask_d2_fp16_w[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21127" *) { vec_data_124_d2[0], vec_data_124_d2[1], vec_data_124_d2[2], vec_data_124_d2[3], vec_data_124_d2[4], vec_data_124_d2[5], vec_data_124_d2[6], vec_data_124_d2[7], vec_data_125_d2[0], vec_data_125_d2[1], vec_data_125_d2[2], vec_data_125_d2[3], vec_data_125_d2[4], vec_data_125_d2[5], vec_data_125_d2[6] };
  assign mask_d2_fp16_w[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21128" *) { vec_data_126_d2[0], vec_data_126_d2[1], vec_data_126_d2[2], vec_data_126_d2[3], vec_data_126_d2[4], vec_data_126_d2[5], vec_data_126_d2[6], vec_data_126_d2[7], vec_data_127_d2[0], vec_data_127_d2[1], vec_data_127_d2[2], vec_data_127_d2[3], vec_data_127_d2[4], vec_data_127_d2[5], vec_data_127_d2[6] };
  assign _09001_ = is_fp16 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21139" *) { mask_d2_fp16_w[127], mask_d2_fp16_w[127], mask_d2_fp16_w[125], mask_d2_fp16_w[125], mask_d2_fp16_w[123], mask_d2_fp16_w[123], mask_d2_fp16_w[121], mask_d2_fp16_w[121], mask_d2_fp16_w[119], mask_d2_fp16_w[119], mask_d2_fp16_w[117], mask_d2_fp16_w[117], mask_d2_fp16_w[115], mask_d2_fp16_w[115], mask_d2_fp16_w[113], mask_d2_fp16_w[113], mask_d2_fp16_w[111], mask_d2_fp16_w[111], mask_d2_fp16_w[109], mask_d2_fp16_w[109], mask_d2_fp16_w[107], mask_d2_fp16_w[107], mask_d2_fp16_w[105], mask_d2_fp16_w[105], mask_d2_fp16_w[103], mask_d2_fp16_w[103], mask_d2_fp16_w[101], mask_d2_fp16_w[101], mask_d2_fp16_w[99], mask_d2_fp16_w[99], mask_d2_fp16_w[97], mask_d2_fp16_w[97], mask_d2_fp16_w[95], mask_d2_fp16_w[95], mask_d2_fp16_w[93], mask_d2_fp16_w[93], mask_d2_fp16_w[91], mask_d2_fp16_w[91], mask_d2_fp16_w[89], mask_d2_fp16_w[89], mask_d2_fp16_w[87], mask_d2_fp16_w[87], mask_d2_fp16_w[85], mask_d2_fp16_w[85], mask_d2_fp16_w[83], mask_d2_fp16_w[83], mask_d2_fp16_w[81], mask_d2_fp16_w[81], mask_d2_fp16_w[79], mask_d2_fp16_w[79], mask_d2_fp16_w[77], mask_d2_fp16_w[77], mask_d2_fp16_w[75], mask_d2_fp16_w[75], mask_d2_fp16_w[73], mask_d2_fp16_w[73], mask_d2_fp16_w[71], mask_d2_fp16_w[71], mask_d2_fp16_w[69], mask_d2_fp16_w[69], mask_d2_fp16_w[67], mask_d2_fp16_w[67], mask_d2_fp16_w[65], mask_d2_fp16_w[65], mask_d2_fp16_w[63], mask_d2_fp16_w[63], mask_d2_fp16_w[61], mask_d2_fp16_w[61], mask_d2_fp16_w[59], mask_d2_fp16_w[59], mask_d2_fp16_w[57], mask_d2_fp16_w[57], mask_d2_fp16_w[55], mask_d2_fp16_w[55], mask_d2_fp16_w[53], mask_d2_fp16_w[53], mask_d2_fp16_w[51], mask_d2_fp16_w[51], mask_d2_fp16_w[49], mask_d2_fp16_w[49], mask_d2_fp16_w[47], mask_d2_fp16_w[47], mask_d2_fp16_w[45], mask_d2_fp16_w[45], mask_d2_fp16_w[43], mask_d2_fp16_w[43], mask_d2_fp16_w[41], mask_d2_fp16_w[41], mask_d2_fp16_w[39], mask_d2_fp16_w[39], mask_d2_fp16_w[37], mask_d2_fp16_w[37], mask_d2_fp16_w[35], mask_d2_fp16_w[35], mask_d2_fp16_w[33], mask_d2_fp16_w[33], mask_d2_fp16_w[31], mask_d2_fp16_w[31], mask_d2_fp16_w[29], mask_d2_fp16_w[29], mask_d2_fp16_w[27], mask_d2_fp16_w[27], mask_d2_fp16_w[25], mask_d2_fp16_w[25], mask_d2_fp16_w[23], mask_d2_fp16_w[23], mask_d2_fp16_w[21], mask_d2_fp16_w[21], mask_d2_fp16_w[19], mask_d2_fp16_w[19], mask_d2_fp16_w[17], mask_d2_fp16_w[17], mask_d2_fp16_w[15], mask_d2_fp16_w[15], mask_d2_fp16_w[13], mask_d2_fp16_w[13], mask_d2_fp16_w[11], mask_d2_fp16_w[11], mask_d2_fp16_w[9], mask_d2_fp16_w[9], mask_d2_fp16_w[7], mask_d2_fp16_w[7], mask_d2_fp16_w[5], mask_d2_fp16_w[5], mask_d2_fp16_w[3], mask_d2_fp16_w[3], mask_d2_fp16_w[1], mask_d2_fp16_w[1] } : { mask_d2_int16_w[127], mask_d2_int16_w[127], mask_d2_int16_w[125], mask_d2_int16_w[125], mask_d2_int16_w[123], mask_d2_int16_w[123], mask_d2_int16_w[121], mask_d2_int16_w[121], mask_d2_int16_w[119], mask_d2_int16_w[119], mask_d2_int16_w[117], mask_d2_int16_w[117], mask_d2_int16_w[115], mask_d2_int16_w[115], mask_d2_int16_w[113], mask_d2_int16_w[113], mask_d2_int16_w[111], mask_d2_int16_w[111], mask_d2_int16_w[109], mask_d2_int16_w[109], mask_d2_int16_w[107], mask_d2_int16_w[107], mask_d2_int16_w[105], mask_d2_int16_w[105], mask_d2_int16_w[103], mask_d2_int16_w[103], mask_d2_int16_w[101], mask_d2_int16_w[101], mask_d2_int16_w[99], mask_d2_int16_w[99], mask_d2_int16_w[97], mask_d2_int16_w[97], mask_d2_int16_w[95], mask_d2_int16_w[95], mask_d2_int16_w[93], mask_d2_int16_w[93], mask_d2_int16_w[91], mask_d2_int16_w[91], mask_d2_int16_w[89], mask_d2_int16_w[89], mask_d2_int16_w[87], mask_d2_int16_w[87], mask_d2_int16_w[85], mask_d2_int16_w[85], mask_d2_int16_w[83], mask_d2_int16_w[83], mask_d2_int16_w[81], mask_d2_int16_w[81], mask_d2_int16_w[79], mask_d2_int16_w[79], mask_d2_int16_w[77], mask_d2_int16_w[77], mask_d2_int16_w[75], mask_d2_int16_w[75], mask_d2_int16_w[73], mask_d2_int16_w[73], mask_d2_int16_w[71], mask_d2_int16_w[71], mask_d2_int16_w[69], mask_d2_int16_w[69], mask_d2_int16_w[67], mask_d2_int16_w[67], mask_d2_int16_w[65], mask_d2_int16_w[65], mask_d2_int16_w[63], mask_d2_int16_w[63], mask_d2_int16_w[61], mask_d2_int16_w[61], mask_d2_int16_w[59], mask_d2_int16_w[59], mask_d2_int16_w[57], mask_d2_int16_w[57], mask_d2_int16_w[55], mask_d2_int16_w[55], mask_d2_int16_w[53], mask_d2_int16_w[53], mask_d2_int16_w[51], mask_d2_int16_w[51], mask_d2_int16_w[49], mask_d2_int16_w[49], mask_d2_int16_w[47], mask_d2_int16_w[47], mask_d2_int16_w[45], mask_d2_int16_w[45], mask_d2_int16_w[43], mask_d2_int16_w[43], mask_d2_int16_w[41], mask_d2_int16_w[41], mask_d2_int16_w[39], mask_d2_int16_w[39], mask_d2_int16_w[37], mask_d2_int16_w[37], mask_d2_int16_w[35], mask_d2_int16_w[35], mask_d2_int16_w[33], mask_d2_int16_w[33], mask_d2_int16_w[31], mask_d2_int16_w[31], mask_d2_int16_w[29], mask_d2_int16_w[29], mask_d2_int16_w[27], mask_d2_int16_w[27], mask_d2_int16_w[25], mask_d2_int16_w[25], mask_d2_int16_w[23], mask_d2_int16_w[23], mask_d2_int16_w[21], mask_d2_int16_w[21], mask_d2_int16_w[19], mask_d2_int16_w[19], mask_d2_int16_w[17], mask_d2_int16_w[17], mask_d2_int16_w[15], mask_d2_int16_w[15], mask_d2_int16_w[13], mask_d2_int16_w[13], mask_d2_int16_w[11], mask_d2_int16_w[11], mask_d2_int16_w[9], mask_d2_int16_w[9], mask_d2_int16_w[7], mask_d2_int16_w[7], mask_d2_int16_w[5], mask_d2_int16_w[5], mask_d2_int16_w[3], mask_d2_int16_w[3], mask_d2_int16_w[1], mask_d2_int16_w[1] };
  assign mask_d2_w = is_int8 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:21139" *) mask_d2_int8_w : _09001_;
  assign input_mask_gated = input_mask_en[8] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_WL_dec.v:966" *) input_mask : 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _00745_[6:0] = vec_sum_127_d1;
  assign { mask_d2_fp16_w[126], mask_d2_fp16_w[124], mask_d2_fp16_w[122], mask_d2_fp16_w[120], mask_d2_fp16_w[118], mask_d2_fp16_w[116], mask_d2_fp16_w[114], mask_d2_fp16_w[112], mask_d2_fp16_w[110], mask_d2_fp16_w[108], mask_d2_fp16_w[106], mask_d2_fp16_w[104], mask_d2_fp16_w[102], mask_d2_fp16_w[100], mask_d2_fp16_w[98], mask_d2_fp16_w[96], mask_d2_fp16_w[94], mask_d2_fp16_w[92], mask_d2_fp16_w[90], mask_d2_fp16_w[88], mask_d2_fp16_w[86], mask_d2_fp16_w[84], mask_d2_fp16_w[82], mask_d2_fp16_w[80], mask_d2_fp16_w[78], mask_d2_fp16_w[76], mask_d2_fp16_w[74], mask_d2_fp16_w[72], mask_d2_fp16_w[70], mask_d2_fp16_w[68], mask_d2_fp16_w[66], mask_d2_fp16_w[64], mask_d2_fp16_w[62], mask_d2_fp16_w[60], mask_d2_fp16_w[58], mask_d2_fp16_w[56], mask_d2_fp16_w[54], mask_d2_fp16_w[52], mask_d2_fp16_w[50], mask_d2_fp16_w[48], mask_d2_fp16_w[46], mask_d2_fp16_w[44], mask_d2_fp16_w[42], mask_d2_fp16_w[40], mask_d2_fp16_w[38], mask_d2_fp16_w[36], mask_d2_fp16_w[34], mask_d2_fp16_w[32], mask_d2_fp16_w[30], mask_d2_fp16_w[28], mask_d2_fp16_w[26], mask_d2_fp16_w[24], mask_d2_fp16_w[22], mask_d2_fp16_w[20], mask_d2_fp16_w[18], mask_d2_fp16_w[16], mask_d2_fp16_w[14], mask_d2_fp16_w[12], mask_d2_fp16_w[10], mask_d2_fp16_w[8], mask_d2_fp16_w[6], mask_d2_fp16_w[4], mask_d2_fp16_w[2], mask_d2_fp16_w[0] } = { mask_d2_fp16_w[127], mask_d2_fp16_w[125], mask_d2_fp16_w[123], mask_d2_fp16_w[121], mask_d2_fp16_w[119], mask_d2_fp16_w[117], mask_d2_fp16_w[115], mask_d2_fp16_w[113], mask_d2_fp16_w[111], mask_d2_fp16_w[109], mask_d2_fp16_w[107], mask_d2_fp16_w[105], mask_d2_fp16_w[103], mask_d2_fp16_w[101], mask_d2_fp16_w[99], mask_d2_fp16_w[97], mask_d2_fp16_w[95], mask_d2_fp16_w[93], mask_d2_fp16_w[91], mask_d2_fp16_w[89], mask_d2_fp16_w[87], mask_d2_fp16_w[85], mask_d2_fp16_w[83], mask_d2_fp16_w[81], mask_d2_fp16_w[79], mask_d2_fp16_w[77], mask_d2_fp16_w[75], mask_d2_fp16_w[73], mask_d2_fp16_w[71], mask_d2_fp16_w[69], mask_d2_fp16_w[67], mask_d2_fp16_w[65], mask_d2_fp16_w[63], mask_d2_fp16_w[61], mask_d2_fp16_w[59], mask_d2_fp16_w[57], mask_d2_fp16_w[55], mask_d2_fp16_w[53], mask_d2_fp16_w[51], mask_d2_fp16_w[49], mask_d2_fp16_w[47], mask_d2_fp16_w[45], mask_d2_fp16_w[43], mask_d2_fp16_w[41], mask_d2_fp16_w[39], mask_d2_fp16_w[37], mask_d2_fp16_w[35], mask_d2_fp16_w[33], mask_d2_fp16_w[31], mask_d2_fp16_w[29], mask_d2_fp16_w[27], mask_d2_fp16_w[25], mask_d2_fp16_w[23], mask_d2_fp16_w[21], mask_d2_fp16_w[19], mask_d2_fp16_w[17], mask_d2_fp16_w[15], mask_d2_fp16_w[13], mask_d2_fp16_w[11], mask_d2_fp16_w[9], mask_d2_fp16_w[7], mask_d2_fp16_w[5], mask_d2_fp16_w[3], mask_d2_fp16_w[1] };
  assign { mask_d2_int16_w[126], mask_d2_int16_w[124], mask_d2_int16_w[122], mask_d2_int16_w[120], mask_d2_int16_w[118], mask_d2_int16_w[116], mask_d2_int16_w[114], mask_d2_int16_w[112], mask_d2_int16_w[110], mask_d2_int16_w[108], mask_d2_int16_w[106], mask_d2_int16_w[104], mask_d2_int16_w[102], mask_d2_int16_w[100], mask_d2_int16_w[98], mask_d2_int16_w[96], mask_d2_int16_w[94], mask_d2_int16_w[92], mask_d2_int16_w[90], mask_d2_int16_w[88], mask_d2_int16_w[86], mask_d2_int16_w[84], mask_d2_int16_w[82], mask_d2_int16_w[80], mask_d2_int16_w[78], mask_d2_int16_w[76], mask_d2_int16_w[74], mask_d2_int16_w[72], mask_d2_int16_w[70], mask_d2_int16_w[68], mask_d2_int16_w[66], mask_d2_int16_w[64], mask_d2_int16_w[62], mask_d2_int16_w[60], mask_d2_int16_w[58], mask_d2_int16_w[56], mask_d2_int16_w[54], mask_d2_int16_w[52], mask_d2_int16_w[50], mask_d2_int16_w[48], mask_d2_int16_w[46], mask_d2_int16_w[44], mask_d2_int16_w[42], mask_d2_int16_w[40], mask_d2_int16_w[38], mask_d2_int16_w[36], mask_d2_int16_w[34], mask_d2_int16_w[32], mask_d2_int16_w[30], mask_d2_int16_w[28], mask_d2_int16_w[26], mask_d2_int16_w[24], mask_d2_int16_w[22], mask_d2_int16_w[20], mask_d2_int16_w[18], mask_d2_int16_w[16], mask_d2_int16_w[14], mask_d2_int16_w[12], mask_d2_int16_w[10], mask_d2_int16_w[8], mask_d2_int16_w[6], mask_d2_int16_w[4], mask_d2_int16_w[2], mask_d2_int16_w[0] } = { mask_d2_int16_w[127], mask_d2_int16_w[125], mask_d2_int16_w[123], mask_d2_int16_w[121], mask_d2_int16_w[119], mask_d2_int16_w[117], mask_d2_int16_w[115], mask_d2_int16_w[113], mask_d2_int16_w[111], mask_d2_int16_w[109], mask_d2_int16_w[107], mask_d2_int16_w[105], mask_d2_int16_w[103], mask_d2_int16_w[101], mask_d2_int16_w[99], mask_d2_int16_w[97], mask_d2_int16_w[95], mask_d2_int16_w[93], mask_d2_int16_w[91], mask_d2_int16_w[89], mask_d2_int16_w[87], mask_d2_int16_w[85], mask_d2_int16_w[83], mask_d2_int16_w[81], mask_d2_int16_w[79], mask_d2_int16_w[77], mask_d2_int16_w[75], mask_d2_int16_w[73], mask_d2_int16_w[71], mask_d2_int16_w[69], mask_d2_int16_w[67], mask_d2_int16_w[65], mask_d2_int16_w[63], mask_d2_int16_w[61], mask_d2_int16_w[59], mask_d2_int16_w[57], mask_d2_int16_w[55], mask_d2_int16_w[53], mask_d2_int16_w[51], mask_d2_int16_w[49], mask_d2_int16_w[47], mask_d2_int16_w[45], mask_d2_int16_w[43], mask_d2_int16_w[41], mask_d2_int16_w[39], mask_d2_int16_w[37], mask_d2_int16_w[35], mask_d2_int16_w[33], mask_d2_int16_w[31], mask_d2_int16_w[29], mask_d2_int16_w[27], mask_d2_int16_w[25], mask_d2_int16_w[23], mask_d2_int16_w[21], mask_d2_int16_w[19], mask_d2_int16_w[17], mask_d2_int16_w[15], mask_d2_int16_w[13], mask_d2_int16_w[11], mask_d2_int16_w[9], mask_d2_int16_w[7], mask_d2_int16_w[5], mask_d2_int16_w[3], mask_d2_int16_w[1] };
  assign output_data0 = vec_data_000_d3;
  assign output_data1 = vec_data_001_d3;
  assign output_data10 = vec_data_010_d3;
  assign output_data100 = vec_data_100_d3;
  assign output_data101 = vec_data_101_d3;
  assign output_data102 = vec_data_102_d3;
  assign output_data103 = vec_data_103_d3;
  assign output_data104 = vec_data_104_d3;
  assign output_data105 = vec_data_105_d3;
  assign output_data106 = vec_data_106_d3;
  assign output_data107 = vec_data_107_d3;
  assign output_data108 = vec_data_108_d3;
  assign output_data109 = vec_data_109_d3;
  assign output_data11 = vec_data_011_d3;
  assign output_data110 = vec_data_110_d3;
  assign output_data111 = vec_data_111_d3;
  assign output_data112 = vec_data_112_d3;
  assign output_data113 = vec_data_113_d3;
  assign output_data114 = vec_data_114_d3;
  assign output_data115 = vec_data_115_d3;
  assign output_data116 = vec_data_116_d3;
  assign output_data117 = vec_data_117_d3;
  assign output_data118 = vec_data_118_d3;
  assign output_data119 = vec_data_119_d3;
  assign output_data12 = vec_data_012_d3;
  assign output_data120 = vec_data_120_d3;
  assign output_data121 = vec_data_121_d3;
  assign output_data122 = vec_data_122_d3;
  assign output_data123 = vec_data_123_d3;
  assign output_data124 = vec_data_124_d3;
  assign output_data125 = vec_data_125_d3;
  assign output_data126 = vec_data_126_d3;
  assign output_data127 = vec_data_127_d3;
  assign output_data13 = vec_data_013_d3;
  assign output_data14 = vec_data_014_d3;
  assign output_data15 = vec_data_015_d3;
  assign output_data16 = vec_data_016_d3;
  assign output_data17 = vec_data_017_d3;
  assign output_data18 = vec_data_018_d3;
  assign output_data19 = vec_data_019_d3;
  assign output_data2 = vec_data_002_d3;
  assign output_data20 = vec_data_020_d3;
  assign output_data21 = vec_data_021_d3;
  assign output_data22 = vec_data_022_d3;
  assign output_data23 = vec_data_023_d3;
  assign output_data24 = vec_data_024_d3;
  assign output_data25 = vec_data_025_d3;
  assign output_data26 = vec_data_026_d3;
  assign output_data27 = vec_data_027_d3;
  assign output_data28 = vec_data_028_d3;
  assign output_data29 = vec_data_029_d3;
  assign output_data3 = vec_data_003_d3;
  assign output_data30 = vec_data_030_d3;
  assign output_data31 = vec_data_031_d3;
  assign output_data32 = vec_data_032_d3;
  assign output_data33 = vec_data_033_d3;
  assign output_data34 = vec_data_034_d3;
  assign output_data35 = vec_data_035_d3;
  assign output_data36 = vec_data_036_d3;
  assign output_data37 = vec_data_037_d3;
  assign output_data38 = vec_data_038_d3;
  assign output_data39 = vec_data_039_d3;
  assign output_data4 = vec_data_004_d3;
  assign output_data40 = vec_data_040_d3;
  assign output_data41 = vec_data_041_d3;
  assign output_data42 = vec_data_042_d3;
  assign output_data43 = vec_data_043_d3;
  assign output_data44 = vec_data_044_d3;
  assign output_data45 = vec_data_045_d3;
  assign output_data46 = vec_data_046_d3;
  assign output_data47 = vec_data_047_d3;
  assign output_data48 = vec_data_048_d3;
  assign output_data49 = vec_data_049_d3;
  assign output_data5 = vec_data_005_d3;
  assign output_data50 = vec_data_050_d3;
  assign output_data51 = vec_data_051_d3;
  assign output_data52 = vec_data_052_d3;
  assign output_data53 = vec_data_053_d3;
  assign output_data54 = vec_data_054_d3;
  assign output_data55 = vec_data_055_d3;
  assign output_data56 = vec_data_056_d3;
  assign output_data57 = vec_data_057_d3;
  assign output_data58 = vec_data_058_d3;
  assign output_data59 = vec_data_059_d3;
  assign output_data6 = vec_data_006_d3;
  assign output_data60 = vec_data_060_d3;
  assign output_data61 = vec_data_061_d3;
  assign output_data62 = vec_data_062_d3;
  assign output_data63 = vec_data_063_d3;
  assign output_data64 = vec_data_064_d3;
  assign output_data65 = vec_data_065_d3;
  assign output_data66 = vec_data_066_d3;
  assign output_data67 = vec_data_067_d3;
  assign output_data68 = vec_data_068_d3;
  assign output_data69 = vec_data_069_d3;
  assign output_data7 = vec_data_007_d3;
  assign output_data70 = vec_data_070_d3;
  assign output_data71 = vec_data_071_d3;
  assign output_data72 = vec_data_072_d3;
  assign output_data73 = vec_data_073_d3;
  assign output_data74 = vec_data_074_d3;
  assign output_data75 = vec_data_075_d3;
  assign output_data76 = vec_data_076_d3;
  assign output_data77 = vec_data_077_d3;
  assign output_data78 = vec_data_078_d3;
  assign output_data79 = vec_data_079_d3;
  assign output_data8 = vec_data_008_d3;
  assign output_data80 = vec_data_080_d3;
  assign output_data81 = vec_data_081_d3;
  assign output_data82 = vec_data_082_d3;
  assign output_data83 = vec_data_083_d3;
  assign output_data84 = vec_data_084_d3;
  assign output_data85 = vec_data_085_d3;
  assign output_data86 = vec_data_086_d3;
  assign output_data87 = vec_data_087_d3;
  assign output_data88 = vec_data_088_d3;
  assign output_data89 = vec_data_089_d3;
  assign output_data9 = vec_data_009_d3;
  assign output_data90 = vec_data_090_d3;
  assign output_data91 = vec_data_091_d3;
  assign output_data92 = vec_data_092_d3;
  assign output_data93 = vec_data_093_d3;
  assign output_data94 = vec_data_094_d3;
  assign output_data95 = vec_data_095_d3;
  assign output_data96 = vec_data_096_d3;
  assign output_data97 = vec_data_097_d3;
  assign output_data98 = vec_data_098_d3;
  assign output_data99 = vec_data_099_d3;
  assign output_mask = mask_d3;
  assign output_pvld = valid_d3;
  assign output_sel = sel_d3;
  assign vec_sum_000 = input_mask_gated[0];
endmodule
