module FP32_ADD_chn_b_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_add.v:352" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:353" *)
  output outsig;
  assign outsig = in_0;
endmodule
